`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bvrv3Ni1R55/fCu1DRsuTUJut7crhUWDHpaiL8Lo+cgH6FHSmzxwfhNNR6NGTUUc
eomoUeqpPd5gJ8lYk5HiapZooNOEXbxqwZN0u92np4xA/qoYxxlrNmwsgmgJd32R
njUWdHTAs8NMMcgiCWceClmp86aj5/Qy8vKj2EvM8fs5F2R/naXacoO+f9ATXGOo
+nXqYhCFogryRImdYLApqvaEWQp+58byCpF4YQm2wAd5iz4A2Uiri+svMdFiWcno
Jf86ibwa5HMIQQlvvjyn1jR6AlgqOqjhXTwnYDY469LmbhoZ9rauQ/6w35Oa2WdA
Hb8Tco0T16U7HqxnLsES7dBRnNgYMaDvrXmorUYtPTMQ2QptEz2JcYz5cMs8TfUF
6S/FIb/4+//W1mp8+9n9YtpYZnsFQxAlZJh9orSSEm8kilyDxEgkuqqw7SgRGju7
DerSSFIVIsQlpoSfl/wtmRW2bDiThzoD+wRvpWOZaRkHsOsjARZiDzWhBIc4SPQm
MrIuC9AoTHOO7vrUjF8eZT1cDpRUi5N6Lk0B4slTtfhXfEKAwafU7UztV0az898/
Cdo1xCuxndxg+53v5PaAJxJ9AwJiekuiWOmw2oL0eEEXRSUKJVwYbe2vFUuEOTI6
tRnWeAb1w8sr8c6jd9zLq9+5ij8ETpRpa0OpK8OkFMsA9+IW6x1UAIFO7oZtknfO
czEP1CVo/y7sG9FZaZllDz941m7AmGiDVychxKoZTzncuNJIMv0G6PukmzaKrFtD
9b+7OP6Q/IZ6kCCkRjANOTbqDNa8G1Eg9uflDiAVolNk2+xe4wRUxcy2Aw8yrPvz
TwVe0pmdbE+SKYv0j9bt84Vpi7xhAe5JhkMxG4TiGoynMG4eHkB/p7nuqNdPhRfR
GxLr8obVzh8jWP0ZOeBNEeB8HYJZjLwTZoTDkmD8K+F31h3bl1OapilHcpSgv3S+
B5q8YsMBpTIiLoteA0b8CPHgwc/mIvLUL5wFsxR4rWSDL71tqk6QOpojY7nWRW6h
8FHFVrfGTf9+IFMRDnAJ2XG70GWHnAtPlwR+V353SV44CchQIYF3LAr74VvhMqme
RKAdC6a1Xw9dNcGcuemg/y8qL44HanAX2oSgwGK/uNQ2rw96l4PZr+J/HZkDC33a
2b7siKfV4KdU9BZgtXdt9IGybdQaYsSe2k/Z2FPBnT/On54L7Ad5gUg1tTdos8Us
S16tGVN6FkSWPMLBP5TpqZsDgoBI3qwVFA4JQ34PtbqnlAjBYnSqzFGAjsIRmjJl
mJrTheomXATijWdN2MWjtrIHQJ4wt52ovkc/5SBqJFU+8ImIDDH8NjgwkRcWAq4L
myh7lIBqRQLMkVHiupvs+2Q7WhynAWTMsJHKGhtyXqw=
`protect END_PROTECTED
