library verilog;
use verilog.vl_types.all;
entity fourteennm_simple_iopll is
    generic(
        NUMBER_OF_COUNTERS: integer := 9;
        NUMBER_OF_VCO_PHASES: integer := 8;
        reference_clock_frequency: string  := "0 ps";
        operation_mode  : string  := "direct";
        vco_frequency   : string  := "0 MHz";
        output_clock_frequency_0: string  := "0 MHz";
        duty_cycle_0    : integer := 50;
        phase_shift_0   : string  := "0 ps";
        clock_name_0    : string  := "";
        clock_name_global_0: string  := "";
        cnt_en_0        : string  := "false";
        output_clock_frequency_1: string  := "0 MHz";
        duty_cycle_1    : integer := 50;
        phase_shift_1   : string  := "0 ps";
        clock_name_1    : string  := "";
        clock_name_global_1: string  := "";
        cnt_en_1        : string  := "false";
        output_clock_frequency_2: string  := "0 MHz";
        duty_cycle_2    : integer := 50;
        phase_shift_2   : string  := "0 ps";
        clock_name_2    : string  := "";
        clock_name_global_2: string  := "";
        cnt_en_2        : string  := "false";
        output_clock_frequency_3: string  := "0 MHz";
        duty_cycle_3    : integer := 50;
        phase_shift_3   : string  := "0 ps";
        clock_name_3    : string  := "";
        clock_name_global_3: string  := "";
        cnt_en_3        : string  := "false";
        output_clock_frequency_4: string  := "0 MHz";
        duty_cycle_4    : integer := 50;
        phase_shift_4   : string  := "0 ps";
        clock_name_4    : string  := "";
        clock_name_global_4: string  := "";
        cnt_en_4        : string  := "false";
        output_clock_frequency_5: string  := "0 MHz";
        duty_cycle_5    : integer := 50;
        phase_shift_5   : string  := "0 ps";
        clock_name_5    : string  := "";
        clock_name_global_5: string  := "";
        cnt_en_5        : string  := "false";
        output_clock_frequency_6: string  := "0 MHz";
        duty_cycle_6    : integer := 50;
        phase_shift_6   : string  := "0 ps";
        clock_name_6    : string  := "";
        clock_name_global_6: string  := "";
        cnt_en_6        : string  := "false";
        output_clock_frequency_7: string  := "0 MHz";
        duty_cycle_7    : integer := 50;
        phase_shift_7   : string  := "0 ps";
        clock_name_7    : string  := "";
        clock_name_global_7: string  := "";
        cnt_en_7        : string  := "false";
        output_clock_frequency_8: string  := "0 MHz";
        duty_cycle_8    : integer := 50;
        phase_shift_8   : string  := "0 ps";
        clock_name_8    : string  := "";
        clock_name_global_8: string  := "";
        cnt_en_8        : string  := "false"
    );
    port(
        refclk          : in     vl_logic_vector(3 downto 0);
        rst_n           : in     vl_logic;
        fbclk_in        : in     vl_logic;
        fblvds_in       : in     vl_logic;
        zdb_in          : in     vl_logic;
        extswitch       : in     vl_logic;
        core_refclk     : in     vl_logic;
        pll_cascade_in  : in     vl_logic;
        phase_en        : in     vl_logic;
        up_dn           : in     vl_logic;
        num_phase_shifts: in     vl_logic;
        cnt_sel         : in     vl_logic_vector(3 downto 0);
        lvds_clk        : out    vl_logic_vector(1 downto 0);
        loaden          : out    vl_logic_vector(1 downto 0);
        clk0_bad        : out    vl_logic;
        clk1_bad        : out    vl_logic;
        clksel          : out    vl_logic;
        extclk_output   : out    vl_logic_vector(1 downto 0);
        fbclk_out       : out    vl_logic;
        vcoph           : out    vl_logic_vector;
        outclk          : out    vl_logic_vector;
        lock            : out    vl_logic
    );
end fourteennm_simple_iopll;
