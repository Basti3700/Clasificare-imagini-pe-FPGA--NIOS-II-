`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6oKFORLk/k+jAjJax2o372zd4uw3CNL/Psd2bcW0XXlHW4o3+n685XjMf6Zh8GLh
2o5Tquwlvi3oTpzCFLwugkw/ksVNYw0Rth61/Lx45UMgmPahNXOEFTbjfEIR1X6a
t2CSgKtAakdhO6KsaeiP/kAHXCXCGEwN/D0kSKr35qdQKM+/IxLTyZNVN4T4zWx7
n85zywMxrtsCOEYhRKx0TFmuKbSD1RxPGHXX36NkIUtGJsAZLAuRfx2RPd7ygkQX
dPCoMFPaQeERTDUfiswtoXGOmcaQqUbvQ+q8lwgc+4GZRWlLutPbu1QiPr6j1l4M
1ZiVgNSFtJiimrQwSxa3+v+P6thzEfNUbT3+7BISC/qaIlu/KUZTmJh9IEc0FePq
avdrYfTK2J5XNSgkCvRlLq+s6IoE8EUIRBSjxf7oAKwQtbk9S+CX6ShpfPRN4muf
41eqt5gds12Bv+ywdXnHJ0dTB5lUeJVeYpsaV6e0KckKKPoBGJ6nbkCbo7Lj7+gc
0NoLOTKRy2mge5+d30wAShGBVqFeA1v8vrJ0deHs14YDFrfq7+W2wzJcJ1LMQhcD
v3LdAOJvEkDSV4jf1KJ178bXMKM3hIY1WR/ZehKKQfGDgkt+nw7jFf5njsCpmC2E
SgKxMq/1c3chHfHqoFQ7mz0kzHIlSONk/T/nw6BbCSdvu++AcCy+zNz/tOZDpzWq
BQUz94mlFlx6tVwQtLmUY+KccV7XubV+SCuTm6cdQsYUi3w4veuWSTg3jbOgRRXF
KZ/OZdMb9lglsvBD/nPMrsoS9eNfWz/4cqMdE9PlA8VCisx6+gfvkubw2THQNTO4
FeRehsAinXiD0sJ8KSaWwfnahju2r2i+JWgQ3TgUMZyEVpY0Hbk6rJgL70ZQrzVu
BzprVjaxmyf4Vwx+S+gfEkCHPd4Afmj4l5KNWXg8Pk83fR72NfWulzAQuZ/YclNI
nROUSGk2UiEP2TMRFDTeFlsoVm1mpghA/TY0fvlEr8Tp5oXTrrfbmSMeL/m1YNqz
Djvgifn1NDKY1swhuEv8OgovBXra3k3MgzcTopuJJ0jGFbO4kgqDrYdji4d1fVFA
92gPLJkyTEpwgHaG450KqZWwLfObqDUmbOyPDyK73EUVucISjcPw7oksOFQUYNC6
OF5Gcaq2ctuArBeqoCrZmHSpERCz9kyfG6bs+wHCjDumJOEfiany8TACTAHfxp4X
58KfhgKXUoE4Ckh7+C6GdxSatYKokyg8YwxHyld5bMj88hha3E6Fwa+abq1doN3K
EyECKpe4ve63EGhyzInHlJabR+HI1wkDemBSIsnoh8tLO9SNClsgd2o8hWASOnUV
MNeJ3+6k4ZcTiOM1Y7MWLeaVejkJ2OJ+yb06be0Mh7ysMQg/dnf4CtgW53Rxtxcs
yZNLSQCtluh1d9JgUzVZYGS2K/8oevPIJFync51xhFKwWrvswzBAd87itv4bpgv6
oJh/dmPuT86iq6cGg5tvRG6pR02VYM1pr5S7vhdGuYYdzAzOGvDtFOysZ7kym+yD
8fi6oyktzjhTGYDiW8UalhfAxH2mYpgdJf+pLAarnDl7Coy/iMOExVjoMZf07PEU
9+a+7L4Cx8aa28OG3A4gFjlDT+L+YEOS+VE/wBYjaUmT0erpuAjqySSvC+SYgBlT
rt7kavVY4xGVjf2FrCxBPxJNuNCUittiLdySocIN9SXZAGCGXr/Q+Z42NAzmsKyL
Xe3L8Kjs+oQKGvemO0N+T/SdQMtWCyQPTvyxwa9h6DBIZMS7ZoULlkJzTyigJLHr
PHLkNuu0b2dRuZ+TNvCaVRrXHjotKPN4lnvIjLVhvf7U1gyQ6/MOieQH4ugQNHAF
ADLGi5eEoGPgUVbfHjBK3EIXJVrYGeRcuYv8hYM6O/qRbMbKstvwcJmUauOxVmlD
HXKZacNsPjg9l9rbtCTcbquWd/EwTRiD7PYpOv7VroN1tik8IoHj6fBloWFyuIcx
tn1epFd5JMyhoYNDAVtZeLlPGjR2PCSkWsb5zCVws+vY2LmVSZVv9fQKoEM5wrzU
hzBjDMAZhejGCAhHV+8U2nFfYrunNlkuBI8b+cPgWsYjrjO/ACU2PkdSKRfWk6kR
3gCSJcuwLhQZD30+M/vXGX3K3ewk5Z+BayaiGozxzIJWti9ePcE2Kc5ZiD4k85l1
T7obectlKpTo0jSEBPHQNzOZOfMKVHaoF1X1zp+zofWR9VZSIjZz2dDOkI6CVNkt
eZS4qDRqAeD2U24ILtLLd2+cUn/zFlZeDMqXvX6B1ZZro0gkAQ3PZxrbMtK4zE4Z
gUAsQ/ws9ssFothK46iqyhvaMHbo/Cd7RKgvG/3k0uNhbqVrqhX4C8WwKkZasMX0
TKxDacxZy5+82CNysEMzrB7zG528F8y950QnPhnMC2+xuaBRG5N3sOryhWI/NG4k
+KDVbEvl55wouoGc7tfcRY4vreqTVPy4ULmUXdvfmgRIrov7cH7+E+AYFY47RO6t
eRQ1NxXi6BeluPC/t35i3csQwbsFP5fNuHHLjAlJzXU4Ul+nT91XKDyN0B6Q8Dx3
bTGaafz7Z+qdWV7mwa71w4TQmF9rZsfGOstlre3Xm3It6mdYei0Jn5vTNgORnEUg
q8IgJz8prWNwukgz46lA5dcAgLeijDCnD2OOwQve96PNYWMBQoEHnS1waRR/aE/5
wyS/fj1CfrTxlWpwuVwIiQWke17GdY8fw1W14xI3wbvAOPra9tJDYHA8uhKmjXi8
8IQTvw0DLGefxBcfdyIJXQAU7lXB79XyEERKdT1cbrbK/ry9L5Ec67LA17ft02sd
AXmHdEhRxmzRRjy6ShRGb45sK9qwp3jXFgNlp7cFLfmoLNXEf1BiKCyeSSkWuRln
Ori+QBI3uKmhNUrLHausqpmearnL7Qd7T7UByipRkUlQMz3bES0634umsHIJfRGs
hGVnxzH5fN7tTKhvfLYw1AFSXtp7rUpBd7OBe0WQLOY6xeTx7jMVPhmFB6UJ+AWC
GApV7LJbXzSQa6pXtKyZ8JPtb2bSVzKcu6rM5UoxwoRJN4lvcCq0UY8UPb0ZJhJe
WXxNHQocAYLadpR9l162nLulnvwh2em/tBLw2aGtkNl53jrTvZtKuEz4OqsCGB3N
xz2UT7t+e9I+KyuRbYbcw3rxeJF+JA54Au/XzzgxwEaKH8knNGUJeR1y1+l5JBm3
LUdgi5FBFqBA8XNxXrISbB9nF7oh2wplZgPpoafWCKM9gOWfdwzGi9rNRarFx2fq
iLgDlYNOvHKr2a2b7imhm0jHBZ5VN57qewXPJdPj8qc9gVvUiMPTQ+x48P76jgKB
9giWvM1XbQxX0nrb2QhXWZ6/p9T/TUpS0b+u7EW5zyaOnrrCDNy7XJ2IREVletDk
7MeLtRweLMFgz1dSD5x/EGuWPEzsCbtpfwRtGCuiz5WJT8xzvLlnh+SNh736blUg
cnacl0oek64Bj+72hP99TMKt5egrRe6XXoN7thGL+vex7UNjPBkXcsOTha0ygkd9
inuagn5uaYLv/cndZSqE6dv7sS+S6agG/Wso3pbCfjiaow7Jw2tRG0L9GvPDaq5y
HZ/gGiNMrNrsGZSXIQbV5NGCgz1ctM8b+OJyU9QnDSFRhJteK+z6hpQHtWnZ6udQ
WMG6jUobzl0bIxT9ZUN2fiPc+i4npMOZBiwRNLWtmQBuEYLghR2HhioSyMo7bo1d
D0pCE6UHtb7+1tmZtw2aIzb16PJECek+UWNcZvG+T/3Jbtfxgj5Z44Uuwikkvx/Y
1uxXYrCicg5KMdC2kc+jnTiLm2tFKVonqmEh8pTDxs7Bb/84fIjRI8EnMJZC83WO
O+gW51ekY1Sb080oLGEwQLcxu5yiRR1KCCfJFePWWiEwQWIQUbIkzo9F48HjuVwT
ouPsawFTWIDbeWYSIP2egKWL3vVupLi2gKYk6oxGtjniqRqTTBE9P79nPaxaalpA
p6VwKNFPFJzj6N+eOKYp5rmJlSY9GUQBOp9FWZCtK+eZH4Ot/l2mjtfTV0Jrw01J
vEeDwveu/zb4BUHHTWwGwIyQP4/TYrzG44FAAz/jDkbxoxUXKZ+qt4CKUtPNiKLm
P3nvoVLss1ehQWWtYTO8MeUYTsyRmr7d97p49f0FGEW1WJWbEU0vidc9F0c38TQ2
Rfqe7W6GvWp08WT751A1KviIqlyEhYZgtU8lSWQjsVoZPlsMOAmklkFeou8VDlIR
5TqUiZHLl5xtIvNrt+Ttvcwm6pBZsX2+MeF6OF+2/eGjaEIpq5DbJp9FrT1DNC+v
WKVKnEZW1oIiwZ0KwJNQMdOGLlXkH79DduZNYKAGZAfX1P+Vlu69kucF+T2SikSQ
PrLgtMQ8xlP+JY6w3dXAAO1JSeGgei/0nS8pVlcpBQ3Ai5Wb5UiPduxhwEaLl84P
`protect END_PROTECTED
