`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fy4p9Q3YRm+XdkkC73bb7EU2a1uec/VOmsJDd/ZhedKFuvmg6dG4eEtEGIu1sayn
h+8EINf+fONdIbswmKTWmz6CICIJiwQ74FJwHld1WR7l6cG56qtHdbOpaApWNAOK
S2z9nuTc4HQMw63Yyu60YOouDArNmI+IBFBbnhqQWcQ+yDtOWB6wAdnnTbK6EDlM
e7X+ZplCyeiqeINWdToQSsZp7ov/0gQMb0W16g0J6ziHJ7joxAh4FziDzqWDxm1S
O/xLzrgFN6aYqySwpGhPj6yGetwusGg1EpfDz4GKcBTIhjn8LvbvWllq0n26TB8n
wnG//01B0ahSbxDNf9sl+eZ62sKNnf8BS7mSwjRRJYSEVyprr4GoQaMITE0C6a7d
96E55AQtWS44UdqdZvUIyHdSWM3ncn/0SBadCd6l61IxBZQtcJw3v0eCSoruJddf
og6OXYiFR1qz+FVC3sjSimJJEc7PHjx7/gBGkwwb7U4fEEMRcBSSKQh156fedfkD
OVZg+NbyCKE7+MokcZEyDHNP2e8YcNTBsA7rJ78AdMbizJpRLuWvOAaxvvcBkxCK
+4txhvu+xon8FjkmJm61SRFm/DAOHELwE+KJkaJT0P0=
`protect END_PROTECTED
