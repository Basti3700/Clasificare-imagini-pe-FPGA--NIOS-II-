`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQINQmUk94Vr0bijaDMvhOLQSS2M1PZEeOmjXGVUfjxvhpO4aNL9fPwt2CEkSHoi
ghz36bJRbPvmI7VQsSg+lzruHXdIcM8C8H9KXjzEp7MM8mi8guzJr3OjbrMOVC8N
6hYjUnZkjMJXG1OpoMPKt7jatthL0VZJLjwU0ZvuuhNQtGJzJ6Uhn53SCE3ac2AH
3LRyUV6RGs80WberRtOdcPWqE+zWTA0z3jp62S2pnmjH8qmR5JIfQBjwchwO+xbk
5Afl31FX0TQcD126WePDt+tkrHCeJeywyTSd5Hubj3l4Ja+/XvPJolTycZ4O8b91
WQkT7ko0Y1jddnpWR2mfhmqoWfMJXcUNZ7T+IOn+s4pXIBvG9eQqc2BHxGaazenO
BVWlqxH4BTy9BlHYe0aYU9LASTsb5woF/Mu15luNo07RYRUkwwsIJw+XLRNxxBmz
KGXhUGVdxVtoldkY3pIbStdytzVCNB1Z3vf4xwg8ck3zHbqtx7O3r3O9bbvF3n70
eICNMXU8EZvbVUuf9ozNrxwVJFg8AEFXVrgHPKlxqX3ScHXjg2DcJEMy0iqlW6hS
CR1q5PggC2Lc8psT5aMhm7OzcfWHH6kaUJqKaYv3xe7zDELRR16owvLviikdtkhe
veWaYvVXlvTXXzvAzyevoBVOsRmlww8fy831ER7dqENHjw1WD8TYVvst2hFgYO0j
brCcawX6Sd1ZKouKODGh1FLT+kT18bTieJZ/KkGNXKBQgU44c88uYBpJB6GyoZ3r
jzjqXSDaBsbO7G9t3Svl45zQeXFKuUfdk3k3iAx0GYIdclToEqxXwbPFxLo6Wlyv
2QXrov3z2nWr+Ok2Nko+4zS5zNP3mnEkIVSqeqioONnRMnPUrXUe8pFAf48drZO/
K58qoNI8WrxgHw5MZY656QrmzIrD9jp56Ugja0115eOWprUNWmw2LgTyX4FUv1Cs
r+HdndJLYQn79IMjTMHPOrgx8rYaYU24N88mFtqdguB6chD6Xk0dI8sHGoNyDU1C
oVRdFCtMSzpLUdLIPNfZgp9TTEvmaWt3IMVWvqJPun50QKSHSO/1INUycHa+trZw
zt//vvrB+Ym8iZMeyMxoWo4YICdOSU7HSmJlrwYptTt7wSJgg9EWmCV+qF9446yO
7agE+/l51LuBq2ao8LvdFNIHZ7OLd1aaiUcPv79OV3R1JrS52rqd4RdQ9mFCGgub
iBwbygTLAM3sxt4taG3VAWeVlD7ztWNHGTmrkP2VaixOpgsxQ4Kn5PSsPT0Q8Tqe
leuxQLA6QbM/V/QQ8HF4jS8AVZhkFQEupj23ewn4dC9S++560kVCtj5Cd6PumKKf
DsJsXsNXQJz+WjrCzGRRU7rqtq49eGDWqO0bUcopc5un3mhZWLUde12cXUgNzYyQ
ReM6kcVLKUucgFZPXxrjt3Z//Uek6jGGowtK28H8Q6WXv9i8fB+jyb+2t8MZ1idn
XEIzitScX0XJNlNIsVz2x92Jt3a41VCkuN98jhctpXJ6sxvMmp+yFLqgEPwjywBw
nqkJsa2VP+e5p51EqxhjA4Ytb9rhFYoT1r8tI1DLUiyh+wLVr4xNS6t2RY/AQQjT
SGG3bV0q3oCNS0Cy/ZP89IAAZVCzA/0IO7UDXvuv1lkPX2PrnNcdKWzzvcQb/mdL
WJXJzwBIGan21mAT3OqwLZLNPQGrXQ7dZ8as3XzR39olBS34BXyoYCJ7dCQuNRtp
rOj+KSj9OjEcuK4KBt03ilppDb4W/5fOTakTmhSeGdg+THp9xKcUaDame6oHWoFE
5+t9Qfq9z/QauulTIsgHVNP7gaKabk8q/R2PkeQO6TLA7G2dVuG1rwVPfCvkIL8T
UjBtiDyzp6gcrTJkLOvUbt5rTLnIKih2G4+8kLtU2CzwYyvLjXn0uGxJQ6a+iZQx
NgLjgc7JKEHizx2xuOOmWvTPWG29PbI98/IhMSgANO5sd/nOLZIyZb04+YVuvwcg
ayvPAYEI+Nm6tZ0C56QeIfO8EkLglP1lnu04pzia15933zeDIOMrm9Cayf2QKl91
iKRW11lqapXzZh2pjgkNqA==
`protect END_PROTECTED
