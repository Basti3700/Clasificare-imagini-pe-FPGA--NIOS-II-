`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rcTA4Q80EEpYCqFiu2bHnbP/VEMGEzhQvJpRMO3A/ggtSLj1cKYaCEyZAYezP8ve
bWIjNWmVpUz8qSehtoIVyw9Tyd0FVZKzGvuBvwZyMuuGlCZUGsQXQn0Nvt106HBn
EWGU525CEHPhqFjq7/PEvhbOi3z6sok3MsoZiPwFSKQ+2qLioKLvCroWBkYm85xl
DcYoNg3ZEetNnaNi4/hJwG83s4ujDmICNcQQLApIiINQ0WgvfCYqVLBLcS3FaNjk
EryUPQoV2iffthuv95E9EQ==
`protect END_PROTECTED
