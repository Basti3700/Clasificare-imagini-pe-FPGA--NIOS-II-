`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRp56Pgl3r6pEw72wnUC++H9SGPBLmrUBf81xG8U1LyKpaYa24TDLVg/Sek1B8Ik
U+GrZibGeEXjs02Vg1wIfvI3opttBsVMY2JUrV5Oz9IDwsaDcLBTQYtfqdiByrVj
KVfdOA0B7WBCTQ6pIetPGDynO9ccfZpI9WBK7eB/uPNxbQJUCm1YmhveDpXlTPHN
1sElFm9OzhLqk2rlEzqOsBupVmxWLo3cIqf7YeXBfb1OneVKFmkVtXCZV997FRt8
/7x0WdemG/9ucF2zqKQDHBvZn9MKtQW6625jYp0Wcg/XMdfrb0/h0zAbXBC2Rq+B
BkKlkejImL3RgjNVXPUmKVpFk2fcBmKmx+wYCbh5nnTSu7jPY01pnmcacM1YF2Dn
h3jOUIutHxAR+tuYFp0ye/bZBIvjFcP6atxO83CZEaXTqH4/oJLTCMIzh7iRV4lf
8rtyPmFGqzhqJUR2Pb4AYK/V4hJ/vhIGBbDV2Cka8OunLKrIPOSMaobEpMjJR04q
M0CGg5I9dPDzlGdjc2zCVfyPhBvh3j7yuBGg9rcU9cFbuyF2YxZM+rDsT3CEzYXQ
Gadi6QGGI8edG93A21A/h/hBc3WBwfla4/8S4WYIz3zcxdHL/iTuJsqCAF00UEvd
Ll2G7Rn8COY4FRjAH7TJUNn3wF3jBgCRWgjaBE0JwrFD8Bo3A4G+nhNk7DYiliPa
ozBJLsWsgeRvyZrAiPNmDTqw5oOCVdwVYt2zNcPgKc3L/l1dlRwlw8zJiwY7IwXl
zuUCyE89h40srzxZ9/t6kbijudNVDYRm5xeMLzlSSiKBZjNEuaLM+1ijx/SvarVu
OgXBBzvpYCojLTkOkAOASA1C9To5xfEOTjmsO8QIfAbBCUWbtN71N2/X2W698U8Z
3sPZTCSeNSksmhnyywQW7T6kVkJXOan/33gYzz5jKCErh3ugyQY5eE8l79Dw1II3
8Y6MyoJcosslGYhebNgiNCrl+Ac3G/S80Mqm7xzxsQWd7CV/uIDt6YPixcd0uuHY
2hotVtNUkrSKdccOfSXOZT5EMrDoqqDo7xuvGPQS6pqHuIHrAVeIpzfdyPeLJi2r
tTCCKNcbKX/Au8NgXWyomJezE2C4yhRiM+JNHgrY/xyWCRbzUBWB4ankxkB444b9
poqYEidccqIUxvWt65HxXLc40ZP7JHruyNsViWm92V08OwIqfVEV7jBDvr7KQIZE
qqMK5YE4YSOovyqaahWaMKhEVBD9bKVsgkekW0d4RQHxdsPYd9uY/gSQxJ+GR0o1
jbjwqHNOGZwWY6QXtyCfa+NYoZZIgr1FwE2YtFuhS0hJl85ip/UvENOIeiPUsdhz
EB+uMdIj80Hc4NAEctB5xD4+LRiZx41g7Cfa7RTmljXHSw+PyiIWeog0k1IkEaBk
bLDxjANN+ndRWBu2K7BE2NFmmYAOwwSnE3b6J3zCrjhF+THKNEJ7MB4/v05DzEDu
eY937wYHp5jfxj0+xnCf4KJSERrBUhrQmBW5TmowPeL3N3mckAM18Zm8K78kGriW
Slwzn3aAVezr/WefaZP1ClxHdaJ8qPVVj/1araJqvmrs6DqVTnjFkjKtNpxe+Vs/
IoCtJQnLDjjnE0vekExEqq1dDV5ZT84yrKA4VNC6vyC1aM1BSrfuc32+CyAJ1B89
HFl/SV58QcSeQaGGB/pEXC1suW+hoKPgYmeX7Fc3A9QJZuxsaD2LvJVQTo1kwgkB
wgqMVdfLUD/1Yj1pzy4oqA8JeIM0USN68SFQFgkuga9jF6X2hBwAuzoJOywbwamC
0CsysbyH2g/h0XFULPnOfQKd3fZRm/bNRPIcb8xfYs/J/xzlTJfvgWVPtsRyIJAO
nmpt264GzpTT9Y0Nu8Fjv/xkqTXf0B3L3vnEqvL/3doOkJpd9IQAKbSDtwSv/LGl
iB6G+P+aDv24rEEHQEh7otCGz7oS1n+IjhZqlqZedsy3881+rqcExzkXc87sjDwL
S9+6RWCxyX1w5/I24iUjsxGEAqkX5IXP52apuxPv/3Tf+oCkZo9JnB8oMw8GKnO1
YS+Sg0z7TEaxoJf6gct9V/mmHS69/O/IHzAZaMEJdzjWBBJ2nCAVRCf3uzGgZ4gb
zCY8BWDWPOED8aJAwVUb+MIZSn9rwS8KFaWeIYa24Xbqi2oJknZ5gVgMTFZ46IDJ
CQIDNWJyj4dwkoxIAha/QBJzsQ07e9biE9gTPJTKI5NDXfcfzewl6oLuNm+a0mfN
33nM/wt6gOmi/mstY9oSNHNdMWloT70odysfk/k3iw68ZUsNNWEfD5s+KHmsH1uT
+oztWSDXwVK0JtyL7ML3ofEK5dhGIp098nn7lSQDnGjCxvvrvzWolPl+DEloqtiy
0teKQkYh6F+J8DrOpt2h8wG5Ex4Q7MgjS8kDcUqc1QiIOuNsJvDgesuDQaW6rsfV
3+n1OM5zuhUImX37xO3hAKsdgOsy7rNyMdP1LBkLWSIKQbw6HJsSnzVKBoOZ5atX
4NzNa1cr0i/M/nX0vnJI+EvYfa07+WrJcvessVe+E0Rxho+K5nUZmhU9KpvRwUPI
R3nO4Pa198CLiz/19cmwZivqwZhVmuhU0RPTk0ioEH885P2MfX8ChVvJ0LaB8NPq
j02x7FWgcWOp0dJz08VDqUDXWEaCxQdPI3NZAFfqCf0BYAnoZDh15ng8g5ZoTvxq
nJnxBtcAtw5i0bXQHjy4zZ99iShC+1zPhvN//UOanikzj3KafbgvMyX2AULyzeia
cmUr8GhqbxAxLJeRZ/S7qQ==
`protect END_PROTECTED
