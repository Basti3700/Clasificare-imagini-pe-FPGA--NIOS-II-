`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TF9alFYBe7k70KvTjK2eD5zqlBghFXLJf4Hyftvf/px+nD8AWKeYQzGg88NrAvQt
YtT95xUXK+HifNw3bn0T7OmCMQyTrZyPSu0DQJJb8mshsqbRKdJHrPgf5Kko/GcB
oRU0o8sQ632HEbiJvD/+KeqcVw8IxdYLdZYzj0BmtLrIEvePEVm3v+ohhfkYtkVS
58OWF5bGlfyVk7Cc+Eed4vqf1RHLGS4XX+xMU4I/q73L1zO9Toow6PxaA7TFJi4V
23+3pa05J9R0oy9LnPFQOZuBrEB/gPcNswFX7siilDR1Iw/S2zg4wE2tdmXnLXLj
OrqxIttZ2CrT4H2hdRPDQ9S56F/fxyuOxCIkYADxZCGEmk0S/EfAEeyKmvpLDXXB
DRoNKPKj28xYlNOaXs+zphDWyPo37p4hJPdW77tCiONU0MepJWlZ/TsSZUBJieqF
zqFq020xr9r/7YnV307qdj1OrvoFwCN7Y/XC8aKuZm8LE2rNoSfknsSsNc0swq+r
0IFArpS/vpml0eR0gxGNQoWoQl8ewbFR2FZNc+dkU0eKUxr2TrIZ4iJJrlVzAwX7
`protect END_PROTECTED
