`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HWuQoi7oa884C/8oA2TDAc1w9j6ljYLU2F099za4zTWu142E6htqHj+vc24xtYb
mp7NR1FfPzDdGrUkzzIhRb1OdGud4+EqLJsPQ2B54deppa1b9kPwSJDLGzb8n3i2
VbuJvC8QIxtEFqFVkfferbvm1J7tdNpA/OfohvsOScp1s9C/vLZjYiBs7cEruNzi
w1AymAzuUJ/OqdUZOwbpaCtR+rfRZAYsyvTvIrR9VxEibZbIYp7GO/FclWR6O3Xx
M1EAAUlzrp5IO11FscwEeZEhbS4hMO2L5K6MN1mCHoPTUHQdAyzHpfV8Ftf0vdzR
/m5ZV4u6Vnyq9SqcvdRUIqMzda521BUT3v19oIxfcVoAq+b75I92HU1A7NanYAta
jTdOwHLWmXEbR4bvYhlVKmpv5p+wre6HC4GMgKzbVdQscBoDYT/MSn+jl9Cm5yIK
QF3oJwmnEetNvW8yODdRQsnRV537JbcRtRE1wWRyX6hY8ZyOh4CYOAKjBvEG/kAi
gTrK9w7lGEqOeyS/Yzxa++dXgWEm1wBw5E+YDjwevc3wILti9sk6sA+zluEPqelk
QtPboXL4wBKqfBkPThqt8OKTha4HQxmOzUjui4HF/eS2I8cd21wwG1DWJKy8G8PZ
mRqzY0A3GKXMYuAttP0dxcruEmpSc5xnhIwJyhVBo0VUXzL6b55lAxIQtQyBvSS+
AAlo2hWCmh2lXRBHFKkWSZZXvBGbL+iq5ZNmjSCDRozXdp7dfm00bd2eb/Fb5Ynt
wOSbRmlh719dc1u99Xe5n8X1kQ5SY/54ikkpJgN6m+9MB8h3TgbatwJZSISAlmRc
C30BMOLjJUugB8xCgRpAnvHc588faqr89skgJQo5GdP95LhZniXp2q+NuTyx2Pcp
vR/F8qxfW9ilkdEbLtkXqRsyuhmtrhrs+RfeHoagqiojBvfrVcV+/IiAokbErAwW
4DyiL77IJYxybcBSq8z4Wc9G1TVPVHWmkTZaIAKK015yWuLubpz/aLTcLy/Bs7Qf
py6t9bNJyXBlKHlKlHeiMg6qCDd/bYyHJUFbba8f3uuhKB2DzDH0yD6FnP9Vm9jD
7+sLT1xscj8HxRUurHnK3jiy5WbUnNRFRkv9585uKFcghYgxH9hZLxnBU5EjfYcI
9mO21Z74DlN+FKXV8gpj09zVWlSEaO5d92ZKNEijzc+HNeDxv5whBETDyh3KszHp
PrzK7u+a91XscCY/GdYPOLL8t1fB5OWpIB66a6FJwlj6wCIkYw0jiHsltG8Qs/DE
uuR9Zip2xWzpOxR3H7g5Sq2qZIbcpfs2fgEcgUjsMjAVvrh/vzpx6MGXudO10L3e
7ScauBaoB7+TYs3xlfe0nTaFzzwe/ex6hd6TXM076vbCrVXKC0moXjfkZQMSqt0c
pd4lNY9eNDaMAoe1WOMsFsMCH+cQf9OgdLi76ma0EqNxgTm0iGlC0PnJ+pROec4v
XqNKqXjY2icImSsEAXpwWduBkaSnu4gO3Q4fsST0DvLoCIS8SCamsEvcnkB29gca
LZFQuM/gT/NswDfT5Q8ihiqrgoKqcdsUfuLojD/ZjkcpZ3Y97P29dOQkWJafbBz/
iVjbrehVKHPngp8k2l1Yp2S9kkgxSvPhQVw1QIPbXZ7GpIX9RdUSQhb7kffMLy07
XoOH9l5TrQ5JkOk1KTMBe8214rcX89cYIyt7gReb/A98Ez+l1sHKrSNOwfQxcNqz
AK2Ip0ZSAqeSrf6NAVOskUp5QSlXY1klj+uwPyCYyY+H0FzXfNNhJOAhDMUYYKA4
I0L/dEgRykQqSY1MNUjYQrNVemdP1WiuMHo2FbRh9p3zAopIKzs0kwoTYtxoQpgY
z+tHeiKQ+uwHkzEeeZh5k+SzBd3hGoVJLgpPCPPRV7rBueOFrShink+20eObmL9s
+PVxVug2dJ831HpNneKc2m/4G7Pfr9Xd42WDMBjHqKqyKWWVf1T0NnbQeMjuvaoT
4PkkOrdV3VdtVGtlUC7kRELxvCKNt2mQ6y1yKZq/5sp02EQllLN6sMwgoydxL+c7
57ZqMq2XHFatflVksEl10QiyPTwZRt3HBoLJ7/+MeMEVMF6i6R3Y3fQCmTp/6yYM
ae9OmGR5xNi2SdsbD/DkanTsmXyaqd74f/nfdX5Lzdi9CwHuIZT/ROkl2ITIpXxR
vhq/2yW/vwnP/eotNBfvUuCLYU9gP6wCWqewgLwrpYqjq2FxuGReUoWtJRNpOjsa
yBA2ITrtLDAtL73WPYFkDPDQT9vfUuyg9DEzsPhvZZYmbSXQ4fGK/JGVok1PQUos
KCX6oKTxDcglia8cq2I/712H3dSTClk0eHLSl5DYQmRIM9qyUw3bij7u3QS7MxyS
MroRZHnndtJ3QsHDouHMhbmv5S2Koyq1ngP398nnAk1y1W5+dAPHppppYb04bpot
1kPQ2w4uX+7z/CmO6bHS5FpR716XQy/nUE+VZ80h8mgnVSEbiLYFudwNUbSBZBrb
EhJDoZluulDptgSp1ZOLVzd+uDDGsgQ/h+76LDFi4GnLVeyIM67WmYQ6HFi1Soza
2i7FPfM4mwRvT5c/yms6cZlLQmQNV01BOkNzXUBK0KcCGBm9q99eTNy2Rd71l+bm
4hlGfi71NHSecMNqe1Kmgh0x3IiUsHtvvRriiSrlQMgsg0Hjcwts8bgRNvaoQ3G+
gSPn9R0pTJO2oqYMyI8E6ypRFjyibfDG/NFgHibiBo6tw0udZyyGYFIRr5JgLnRu
ZW/nXiVSvGZ62PSdGY3WBJYxLFBe/7H7UAlVExNdSpsRnfyTx7BnpG+E/oq64a8Y
01opMxRzYM5RAyhNuGVhaTe1NOzag2ubm3pS2qsDA5qBxlhTqU3NaBuabI9bga7D
tnuIyhCnyQWRAW97XQtvwFzhhpi16nIxJgjrYh+t9zk8DH8MZp4y/qlZyeQymJah
o2yj0JzCSJl07vcJK/R+fZBsuZwQg5DDkdv5q6G0aN9ewcajxuqoi1/vueaUNtV8
F/BZlXAzXfcoQYdT9yky2apHJOzOQyzeiWzxyYurC1GgObNaCo+bYcRchhlcf3RV
NHLYG6vPjk2YTItYiN+zzls7wc/qGjggcGaLyRhkOsOvK+h/vNh6ZN1aHRgFdxH1
Tkx54H3n2b8U4oGMjWnVYF8CUxjSZifjBomn7DVD4zM8u7LNz5/6kdnruIbMvwDY
Re66IBuRlZM2ARr8tw/HubifgyHmdjreRA6GZ53Ebv9Mb7gLmnXKE2SThsPVnMDi
+a6Ip5TfT+QdgMNU29XZN1j7UUze9Xy8cMCLrNuQCLht4rOkZ4ScCsVernRwd2O4
sBtc5ORKF8tPaPcaUG3vDPolTdkQIQSd7U6X2beIY1/d6qoJJN3Vqoy+kmaUToR9
fSsvCM0XkLD5B83Ng71ymAp5m6w4fP1BFxsTgpC8dqAjVTQHS58ccobn8rdlA/Qf
My/ZxBrRnGgfEJ8xpF7KK/ckWn3NKRNw9QoeIm6sIWUxeb+iDXXshW/iISxH2pag
X5eV2NxJpFsUG60Mljmwz4tsRnEWRqVtdvbm3FJU2lGq9RN0AMn+VfU2Wf0TB8FS
mM3ZgvN94ib6//sRJo1Yx/SLuywBrvi/0kHLZ+HTy2LEwYCFDMlfxnBpg1wYIN1f
5HFDrSZdtBDVaNOWVAqyQKlzdaiSI+G1TcDtfRd5yMMGKPde0080gDeqZWFo5sWw
LZLd6kMJixOkpcrV2ptHjzOxg2zHwYKzxd57U1Umokniqsm2pJgBQ8Hgx1kVyQqy
2QkAXpTZeQcDESEERGirs86+8GliP4IFeQ1CCd0SqIqS4xUi+cvLeIhig1o5AFe2
AEYeIjEnOnl0juhx9Uc9s6LEjW6PYObORBk/XOGnrm45vPa73FqqB4TH4pH+u8yb
SGana67BpB2RuUG/WPEZ4AhFDzLbVZIhMt6tCqDxc86035daL1BtqPgNTOG5oXnU
IpzHpYCDjZXAJ3mQwQT87FpA/8xE0fU2i7HNWJduxPgqh+rMbOE62olDZKaAuDlX
4eG/C0vK/yp+a7+nF4FyVO/GRoZ2uILXnBjLoWGJ+H6HWSXYugG/tTFJlpPvl73x
xnnMOZoixsBHsfZ8qqEQT4e8xVirJPl+8lpC0rK9d52F2aCcSFPyMa4GRyhNiERk
kYdeMHSv/fk8MkzU9+y58GGV0156cXxMnPrszGTkrLJ+tb+YCNVsQshd0NiGCBtK
/6dWcxWf7QnhEdW5vJb25Q+aPIrZLZAeQZxdGyPeDAzRH5dbCUGmz22KF3A5ogsT
ouemdXzfVcUT7YuacAYj4B+3RKcqgl9ycsbjj7UDIeHVXj8XJH6ism8YD8MMX7om
W13vAZeHBk9vsKH1xSSvHcYfmArsFDdy7+r7Q+yi7rAHZqcm3B4JIXX73YmKadPq
SArzQ21RK3MCygHTBSLJzKYIWx5jTH9JvrdcAF8+nAuF9/w+0IF7RHzLHkMiCOey
u0uBToVbM96bcsx4gcLFM+EHDnTGH95ryTq+Tw3fsF/16juA7auWnOY3k/iitvSr
FJPj7MkIIdVGP42xu5BR/Ndc2G87OQhuz+6itC1Xsl0MIqGruxT6aRB3eslIDIKV
LS6tsfUIKTSao9WfX27o6YJFYpun97Nr2v8y+ffnRBhUVDoa+YOpwfeyLEcovOOY
N33dP8TnhcA2/yB1ty+ej8AQS/nVqkdGSGAlg/sqSRLqxv9dKVzqDOBcQkpjKZ6X
mA2qzh6ty9QMjCNQK/CQDiMSk1Rqj5REnEDZxK9UNVPGyI9sLMqd3cpXqv83bPlB
dMG36VFhLJmDIhVYPArvXrf8HxccDzFIqj4kD7ABAYjsHTNCtcfj+TEhr5Uv5hOg
9Bg/3txSZ/qwr8PlfCVt3dKRMfaU7w4gx2Icb4Hmh7A3/0XSRLCa8+UIydhMQFdJ
1tqc3cTqobSFOwk54vRtBDOsK+BMzmlZXoKdq3XU0uydufw1GGr5fMYvjmttN+cy
AGx2QNXWmouRai8RRd/E3nJQhzi7X4vzndcRfv6tmMMGSCmS3pHu6oPp46OIMmx3
FErk3a5UEfDPg/VeIPoUHfzctPk13vFtJb2RPnilKCUJmGOmswNbIgSpVlO/rM7m
CTFC4ze1eNsDhCaiVT/UR10cayFUMuAJhRjr7RYzWS+kMdDU6oCrrelMOG2Cm8xi
26VM6N4UhVtzvHUutLHSLDF7DAlJ0WM7XeaLQDv9gsoLCd6BTu+vA5kcqo76QEGj
Hfwi0rmfyU2D107vcnqZOizcynJ3ofFXaHt2ARrqjAu8c19n3I71uqurGH6sNUGs
GyCLsCP7XCY7PvTiZxcYFaE9+OBnA9wvROi+eVvbgTtM4JRfAGOh33Pkbu1/8LH9
XVHkJMP8Gl8dIUzJN3rISGRo4LvaUAlPs4AXa+tvLMv1bipbAVTht0ncBCiNh037
ADf85pCiXCn7Rk22OZyRMMTDkkuU/gYuZPoJgr0s4W6dUAFIWhRRn2Hv63qi1BsC
HE2XO4/qJFYfQr4A2NyN2qYvSqcXYzUntCtpUClWUZBsj1ZXqSXgRPrvjSKxQyMB
wN48d5wO7bvOAcoYPWOB6KtEpeyze8aagT97YArbORt8Jwtz8irrqRSoXR50j80A
b6hjSf/mdBa1VP4VGf2zIo/EUj/n64NcR3XdA6euypJ8zG3dmgvojm+Iu1Y+rYGS
PCmY825TI1ouWdmE61WFTeWxD5WWWKIf4WiCQ6UETm4U/m+zWActdLbzc2S4xeuk
khJBHXXOF33vrBJ1U+ZL9cGp4fXBqJPsCWupD6xkeKviZL5rv86CG4kq7IPyVcjI
eUbyacKsyR5sCkv3dutqqC54WgUZUV6EWj0pNVjK3bKjW5nqobHV2T1XYdkPVMwu
Gre5vIOrl2DfKuwfbuBiKHTlpAaCWppoJGM9ExIHCrjgzIhG6o+EKWK+nEc3REN8
jbEmxkUsi0VdrxJTWeA8stZoBGLvYr9gVW+nCaJHevn/jYOHMnH9iTVALy4+a07O
y2fE74Vbag6Nw+wpvqsFtfruOtUSQF3141/FU3h1WZb0W4Z4xjD6Xtu653u7nNgt
hHykq7D6mZw/mTaKPKWk22v/MnNdmG3+XPHtUvfLMKhTMAxECr+BICS237vtoalg
NazYBlk9ODLjGeLwNtBnQYjsrQpGa27TWFg9aEBQm1mDSoVI5Ff+iVz0WBm/FVGq
TodsMyPALAeCfyF0UuxG0TwSEDnhJbhJrE84l+kfTF4iuHZeWBgCd4Bpux37TDtm
wag5TdWHx7qGJ64lMNXQkv9szRKZPg3OIZmuFYPFe2PVM6GQIG3WHuTa3OWKs04C
r+f/6LRBeT8QMpbDvzZ/zfLG57XDzMAVkMSvZnfM3gdzlYE1oH2GQ95KOQfZ9m3A
6FMVKRiIGAONWluiu2svkhBXXxQGM5Je010tPOF4+msHXOreHGuyUNv6UZJVJjbG
08n2RDMKZYcgpJytLiJ/rG/UGLFuugjvZ2UzOxJOPzSAk7q31OfAQzk8h6epR/6y
BKSENA6PpKOKz9rLDPXYIEAZhFZtHFdU5EXrkZAPMLRo21QQ5C5GGjHxXDQz/4dh
UO4RgKG1XIyIX+RtsbfKn/FZ8HWCWtbU/BaGmybxs/W6ULSCY2Gg4J64E71ku9JS
Antj1N+yqovuF12X2dTGbGjAWn7SWoFmyW3Q/cHyGHytauuYwYj9TbcVjn+xE6s0
6TQGTaJ8Eb908NGMGvYPAcwlLnCnOpk9tD9QkXz1JlM=
`protect END_PROTECTED
