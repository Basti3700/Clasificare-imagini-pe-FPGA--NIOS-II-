`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XDQR8MC4OeVh8K1ZcKvGrzAEk1bJFsHu8bmSkKqIhF2BjR3z+DTJJndh3YiZoBLw
PkfG2J1m1XlmdVT0Jg2uc7Om3lPp7w2ogNdPzCk186XJuTP4Rbkl52F6LAQzOlL6
RX6d96VsMQedgBrJ1oLknqhlUvuUXwKyHcPzUkD8mMKZghsCFDkeIWbWwtIvcvSI
w4I3VsMmJLOYZaSLWnGKsnchA/Krt7zqrCnrF1SvJ7IoRmLzAgNnLfZ220znCsAS
G47sKKmMgeM41ll5r6871mjaDVGVB4CDDL0L+EL7KD+kHo99VO6JiR+jdcp1pkGC
/IG6ZMOuNE1VXSdpmGQ1osbUrXuAq8wO2Y62yOwj/evJDxgr2oebaU5BEzJlnLVj
gXQL3XISttJPuUPUTujYPxpGAvb9jnXaN+rohmtc5fKh01KHd41JWHpwMPfNm8Vf
cPtiAzTJqNRzhTLHy8Dm0PlJfzQ1zt5XvIWcb5CD9060CaBMbzv2dXzji+MumuYX
eYGPUbg9S7aDz3XghKEhKHLcLHpDlblJhv9YoTIqUqAFyueds639qW5GnXHlMyV4
8dOMOZ9jibl5EF91KU2bH524CDmO97kvlTJ0/MB4vbvhh/QljqnU37Y7hnucaIFQ
bk+iVQ6miJWXiMB38+3jjw==
`protect END_PROTECTED
