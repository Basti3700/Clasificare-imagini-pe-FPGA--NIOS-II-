`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2z5o7y89ZifpIhc4y/OXKwT3MBriUurpevxaBEZFJGBQrDwBFgX30eU2sqwESfR4
zqe4k4UZ/jaZbwwwd4si7z76nskvBzy9Wfvx4emI2dHUl5Ix0635RGueK2Lrjb3M
ZfoAwqypBlN+WU9zqYtNpHIty3R3OP7rbQGPd20dOC2wHh7lrbWkDQ1HzF495Ea6
mtHrHsaTrscRZe9FIUUFcBJmbTII+Df1OCdwPhB3XvyMTDV+yBxei2oqov0rBEBe
fiWAeDQeLsJOBhIKaCuK+gZvWiJoW3NdQJm5IZKLwovrryoOoGitL27KEK7q4eg0
JbuoZ+mWFJAdcbosnqfc7h9jmWJAywNbRMb92K84P37N7vwX+YWg+UQQ+UVX9XnR
YnQAsGJYGUwmi+ggZ79sEFbRrHcq6bIx3mXyTxrshfNjIxSRbuByCDCLsyT2i+/N
AzSm8ubtMEOORcD8YFGI3CQ6yXu+2WGNa8NH8xTKCMm0mc+vYJHSPTaBpgfn/a0t
GiBjd4Zl5J8ZPU35g3I9HnFu+jaPOffaDFVxy1uU24ghM9jwEOOfFEg8ixPB1+KC
c0s1W3rJimYJufgOWhwRGbjzbwh6bLWJICS2Rcry7ByQpF3VMeu2TeABeEr+M1S8
ovXbdhSPDDXIoKcgWtOAfwZuMH2n7+zXV2G6JKHmN/Xb/ErztSpS/jZXERv8jiC/
2bQDPl+kaL+HRsTB9JqGD+Cr+SUOMi36x8oMvGHTD6Qs2VdRT33ibRwxkh+HuKC0
/MeY5RdULocpI6KyQnWOWhGhC4xgVGp+4waEXYwPZ9pF0cn371630qxrwMO/qS89
J0i2TY0itqSiIcUvEKitCUonEY3A0LUzV/cBPOm0xZi27SzSuhu2LATqNMgszt6i
l4/tenNfpSGQuaekLh2aBJCgV9eUePjlqQuD4zyuxEQ6uLKPy2lU0v9LvcpKMUK2
yBJ6MrMVDwsgXHhgGIZxwQCIGFtXcFsPTSNkUsqUSgdlfziLj4Iy1lQYj6F+HdMV
WnLcgOOhYwoxtMrME5d8aJWsYt83vPRQ8odnJTL5MbjZuFJWzFFiGnqrH6fNezkj
E7LtKqlQStXASLylIiudFO0azUecST5iKPaQFQKfhZ+4zH+U2DWMvOk8JNwHSg4H
S6pcP/IDiiXJse69ExbZIiYhrD/ZvkGML3eERcuunWEBCX6852ymJFGfwbTA5ARO
RsyVO0km2HCg1fanuR4kTUKAqnsAxPHA3DSP8SWvQrJLJ0S6AhyxDzxoCHHNhV/9
htt02MPgFUfGCQAfkwiexkRXME9xpgslNisqbVax50DVXLHgKwH7YtsTRiSRKnfX
Q26ozWBptNatOlinGU62Q5/e+lxhAH3x1YVYwrqnEKcWjE8CNRDGL6xwm536rhah
cOXNQEc8Jvybr7eHqkKa9xqAyhfuxBjunnPeKJ7SYwaH6FLtwKEv31mFtqEyeLVY
zqTvW1oLIqje211JLV+i9G4/GOEAHKGVanm0QVtla06zeSdl41JQpi7tmksxqy7Z
9Yw5vURSlzrRoDPN0Z569F4nEUDgLJG2ODKmvGktwFCzLYoBZrwZaDbFNBSnN56z
3O4f+BUcuKbd8N4gKLusyS8+sKlrlODplzZxoc+2JGlmgpUCb/6mh2DM3RsxT0/h
KIZmU+VaG0Uie1AVZiVFyBy1SsBQ3JtHLVgCv/gBX9rzmta6F9m7e6WkwdvC0cX7
/M3qiFjPepQe1V9mb8ZeIfCNaC4N37P+4I5xWwwQkRmjTKGQx9PENXN3Vh9xlk4A
RocrVIdrS69w68JrAUy0O6q1lT+qZlW4Nszk73n6o2xpf/MJCHYOCl/zmtWWcEUC
ttKZ+KU/dR+4woUR0u/J2g7JrQde9OlkXEvur4FthpL5F3xDYw3ocqk2i8P5q+NY
/ezJhoGPSBeLtvqS5XXbjxU61mxo3Je8v1t2kBdzW/O2nYFp8ZNjGa8XyIPzGKTc
W75kiZlwSKQHCLxZE3uT3wDfgtX+sOu/Sb8D6jiB1TQCFb0vAQaR5rRA2SfGj/TN
uRddBboh0AKFWM0XfAFlFHfMzEtUUQpXJwxUDZOmxm0tAZgMG9RegMMLpkgSX3ct
PAyOBE5kAlSosxBA/F9Gf0THeu8x1rpI6mA8lxctHJK+nwYgxkpdGncib6NyTBtH
eraeeiHAFOfEDwcBKwxa0HJIekEBg6s6P9Q0dBRS39xNA2vYHdC5U10WrV12HF1i
N79fw0uyv2N28Ay6WXsirx8rE2nQ20OXKj3tOWHUkuQHD8e51YCgrQ8rspbgXTHe
rULwgOYtlOSsETvqnNWb4GsR1P8ht79gWpnvuzcFcQBwZ7fAVF01AZ1fCijh8qx7
hT0NFg2GCNArn1xcDC7P8/l61NTsiQQmYk5dpvF5ElYYZWd/uuG0Ap5R4sBlnqZP
BECyKrgLGSSQyp5DubcumzosdcmCaMXcMrHFP5d4UlzNieCPZtz8G5P/5Klum493
V2ekcy5+Bsk+Oc+Jz7ijdUQSUUcJTt9+Mlqa9ODEDXxlaJbMUBZ6dbZA3CHvxIw8
34rHVMYZCTABbusH8XPQa+g0gXXfFkkNnlQh43o2a6oGFIwOjcHfGPJViRXaIQMd
86FR8utZKviGaxCnp7M/e5wqT4b/Yfii8OQyE3KVMWc5yM/zB39whbWY3cx4Zz7c
wOwMc3gduZHBx5h5ETFebY4GSmcDTdzfjnGrc40d5tImi/iavnUA5ZHEFb6LEzn9
jcUhX6I8yn18g0AbNEgap5/kbTWJH9jxVCEGX4g1d9B9Z47RgBsFq0fEIJmfUg4i
rGDlkcbK95ScEZ1EKa37ZmZAKDzqFxPUXCVwyD2pd+72/HueLe8bE568exkCJ9pW
YR+d71Q4axrHQT/l9z89UQlNJD4kCRpftRUxCqjxZOerqlt9XovmmGFchE2M9wRg
i5NEZdgyumNM2nLNAWHEZKM5YT644rPsR60cIxUEshhyuYVejONJ1OwQTS8c6Rkd
4xhWjBZajD7e27qm/Q3bPXHcRpG1G65HDpq8fOi0rWf5xoky+UUISVB7XF6+6EfT
ExX56q3igrojvcQzmfn+zBoYn/6l2tkz+bAMU/sljqTYC9dh3Adl8rpKBi6Ix15A
rxeXWIvziuMxoM1gpVvb73ydUvUGAFvvvF6hbjXYbTf11R/md0AmzCtkmDp/GrmZ
0d2rKFKDK0csiVlhukX6QAtRyB2i9OhJKFOAAzbIOFb995MP7O/o4dvdtEKNDBeW
dHJ29S5ufODc6GQ9YDKNgNaIG1kiG7EgB3AC/GWOlUAa0LV/idzQVuzZH4iE6F8j
eBSjj17ksSpd1KVnbD7pxb7u7PUDsj8uYHTAZSsLW/ECsx/A6zBC7s30+5D0kByF
8hDrFiAAusD9f1zTeMRjXsRhwquJlyk8I+Gm/0tTDabzIYKgpp2i7e+JbnnHPsqU
o6A7jEq7eQKjPmT3VKQkuzUAVvaAKaEj9ZGFitQ37SkiWI8AhmTg16lWH7lTz9u5
6Dh6JDgoZ8sUT8K7t1kjLO8f0nfR0LwPwarRQv2tu8MoqPRgBjtbFdhTC+sb1eaG
RaLWV5CSUGe438iw03rIXKOKesEy+RR1oXWFaOlrC5kVG8Hm0PX6ZVJoh7KFRHEJ
EY4nNbPHWjD0lnUuwPzYROO0nz02S11WxolZ8gOke3Yz/BSPo5t6DDTqg2guj8RT
vPnYy6oTeUTAsLrMthOiWXjeJ0uTas3T51Kr6vs+SaAhlRZS9939zonVIuzh+v/+
IWekwpnFGnK5VlquidZ/dfQ/dfnKEYXddmPMZL3jKJmkPK7wL4enzj1XeNMFvwYc
SfzZXrxIG1/yhSnekd0OuV4bYpDyCZee8jZnQBenLD+Kpsg48sy5Oo/RUqtrAfCI
OrdXpZH8zw+MA6c11+D0bA==
`protect END_PROTECTED
