library verilog;
use verilog.vl_types.all;
entity altera_pll is
    generic(
        reference_clock_frequency: string  := "0 ps";
        fractional_vco_multiplier: string  := "false";
        pll_type        : string  := "General";
        pll_subtype     : string  := "General";
        number_of_clocks: integer := 1;
        operation_mode  : string  := "internal feedback";
        deserialization_factor: integer := 4;
        data_rate       : integer := 0;
        sim_additional_refclk_cycles_to_lock: integer := 0;
        output_clock_frequency0: string  := "0 ps";
        phase_shift0    : string  := "0 ps";
        duty_cycle0     : integer := 50;
        output_clock_frequency1: string  := "0 ps";
        phase_shift1    : string  := "0 ps";
        duty_cycle1     : integer := 50;
        output_clock_frequency2: string  := "0 ps";
        phase_shift2    : string  := "0 ps";
        duty_cycle2     : integer := 50;
        output_clock_frequency3: string  := "0 ps";
        phase_shift3    : string  := "0 ps";
        duty_cycle3     : integer := 50;
        output_clock_frequency4: string  := "0 ps";
        phase_shift4    : string  := "0 ps";
        duty_cycle4     : integer := 50;
        output_clock_frequency5: string  := "0 ps";
        phase_shift5    : string  := "0 ps";
        duty_cycle5     : integer := 50;
        output_clock_frequency6: string  := "0 ps";
        phase_shift6    : string  := "0 ps";
        duty_cycle6     : integer := 50;
        output_clock_frequency7: string  := "0 ps";
        phase_shift7    : string  := "0 ps";
        duty_cycle7     : integer := 50;
        output_clock_frequency8: string  := "0 ps";
        phase_shift8    : string  := "0 ps";
        duty_cycle8     : integer := 50;
        output_clock_frequency9: string  := "0 ps";
        phase_shift9    : string  := "0 ps";
        duty_cycle9     : integer := 50;
        output_clock_frequency10: string  := "0 ps";
        phase_shift10   : string  := "0 ps";
        duty_cycle10    : integer := 50;
        output_clock_frequency11: string  := "0 ps";
        phase_shift11   : string  := "0 ps";
        duty_cycle11    : integer := 50;
        output_clock_frequency12: string  := "0 ps";
        phase_shift12   : string  := "0 ps";
        duty_cycle12    : integer := 50;
        output_clock_frequency13: string  := "0 ps";
        phase_shift13   : string  := "0 ps";
        duty_cycle13    : integer := 50;
        output_clock_frequency14: string  := "0 ps";
        phase_shift14   : string  := "0 ps";
        duty_cycle14    : integer := 50;
        output_clock_frequency15: string  := "0 ps";
        phase_shift15   : string  := "0 ps";
        duty_cycle15    : integer := 50;
        output_clock_frequency16: string  := "0 ps";
        phase_shift16   : string  := "0 ps";
        duty_cycle16    : integer := 50;
        output_clock_frequency17: string  := "0 ps";
        phase_shift17   : string  := "0 ps";
        duty_cycle17    : integer := 50;
        clock_name_0    : string  := "";
        clock_name_1    : string  := "";
        clock_name_2    : string  := "";
        clock_name_3    : string  := "";
        clock_name_4    : string  := "";
        clock_name_5    : string  := "";
        clock_name_6    : string  := "";
        clock_name_7    : string  := "";
        clock_name_8    : string  := "";
        clock_name_global_0: string  := "false";
        clock_name_global_1: string  := "false";
        clock_name_global_2: string  := "false";
        clock_name_global_3: string  := "false";
        clock_name_global_4: string  := "false";
        clock_name_global_5: string  := "false";
        clock_name_global_6: string  := "false";
        clock_name_global_7: string  := "false";
        clock_name_global_8: string  := "false";
        m_cnt_hi_div    : integer := 1;
        m_cnt_lo_div    : integer := 1;
        m_cnt_bypass_en : string  := "false";
        m_cnt_odd_div_duty_en: string  := "false";
        n_cnt_hi_div    : integer := 1;
        n_cnt_lo_div    : integer := 1;
        n_cnt_bypass_en : string  := "false";
        n_cnt_odd_div_duty_en: string  := "false";
        c_cnt_hi_div0   : integer := 1;
        c_cnt_lo_div0   : integer := 1;
        c_cnt_bypass_en0: string  := "false";
        c_cnt_in_src0   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en0: string  := "false";
        c_cnt_prst0     : integer := 1;
        c_cnt_ph_mux_prst0: integer := 0;
        c_cnt_hi_div1   : integer := 1;
        c_cnt_lo_div1   : integer := 1;
        c_cnt_bypass_en1: string  := "false";
        c_cnt_in_src1   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en1: string  := "false";
        c_cnt_prst1     : integer := 1;
        c_cnt_ph_mux_prst1: integer := 0;
        c_cnt_hi_div2   : integer := 1;
        c_cnt_lo_div2   : integer := 1;
        c_cnt_bypass_en2: string  := "false";
        c_cnt_in_src2   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en2: string  := "false";
        c_cnt_prst2     : integer := 1;
        c_cnt_ph_mux_prst2: integer := 0;
        c_cnt_hi_div3   : integer := 1;
        c_cnt_lo_div3   : integer := 1;
        c_cnt_bypass_en3: string  := "false";
        c_cnt_in_src3   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en3: string  := "false";
        c_cnt_prst3     : integer := 1;
        c_cnt_ph_mux_prst3: integer := 0;
        c_cnt_hi_div4   : integer := 1;
        c_cnt_lo_div4   : integer := 1;
        c_cnt_bypass_en4: string  := "false";
        c_cnt_in_src4   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en4: string  := "false";
        c_cnt_prst4     : integer := 1;
        c_cnt_ph_mux_prst4: integer := 0;
        c_cnt_hi_div5   : integer := 1;
        c_cnt_lo_div5   : integer := 1;
        c_cnt_bypass_en5: string  := "false";
        c_cnt_in_src5   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en5: string  := "false";
        c_cnt_prst5     : integer := 1;
        c_cnt_ph_mux_prst5: integer := 0;
        c_cnt_hi_div6   : integer := 1;
        c_cnt_lo_div6   : integer := 1;
        c_cnt_bypass_en6: string  := "false";
        c_cnt_in_src6   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en6: string  := "false";
        c_cnt_prst6     : integer := 1;
        c_cnt_ph_mux_prst6: integer := 0;
        c_cnt_hi_div7   : integer := 1;
        c_cnt_lo_div7   : integer := 1;
        c_cnt_bypass_en7: string  := "false";
        c_cnt_in_src7   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en7: string  := "false";
        c_cnt_prst7     : integer := 1;
        c_cnt_ph_mux_prst7: integer := 0;
        c_cnt_hi_div8   : integer := 1;
        c_cnt_lo_div8   : integer := 1;
        c_cnt_bypass_en8: string  := "false";
        c_cnt_in_src8   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en8: string  := "false";
        c_cnt_prst8     : integer := 1;
        c_cnt_ph_mux_prst8: integer := 0;
        c_cnt_hi_div9   : integer := 1;
        c_cnt_lo_div9   : integer := 1;
        c_cnt_bypass_en9: string  := "false";
        c_cnt_in_src9   : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en9: string  := "false";
        c_cnt_prst9     : integer := 1;
        c_cnt_ph_mux_prst9: integer := 0;
        c_cnt_hi_div10  : integer := 1;
        c_cnt_lo_div10  : integer := 1;
        c_cnt_bypass_en10: string  := "false";
        c_cnt_in_src10  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en10: string  := "false";
        c_cnt_prst10    : integer := 1;
        c_cnt_ph_mux_prst10: integer := 0;
        c_cnt_hi_div11  : integer := 1;
        c_cnt_lo_div11  : integer := 1;
        c_cnt_bypass_en11: string  := "false";
        c_cnt_in_src11  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en11: string  := "false";
        c_cnt_prst11    : integer := 1;
        c_cnt_ph_mux_prst11: integer := 0;
        c_cnt_hi_div12  : integer := 1;
        c_cnt_lo_div12  : integer := 1;
        c_cnt_bypass_en12: string  := "false";
        c_cnt_in_src12  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en12: string  := "false";
        c_cnt_prst12    : integer := 1;
        c_cnt_ph_mux_prst12: integer := 0;
        c_cnt_hi_div13  : integer := 1;
        c_cnt_lo_div13  : integer := 1;
        c_cnt_bypass_en13: string  := "false";
        c_cnt_in_src13  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en13: string  := "false";
        c_cnt_prst13    : integer := 1;
        c_cnt_ph_mux_prst13: integer := 0;
        c_cnt_hi_div14  : integer := 1;
        c_cnt_lo_div14  : integer := 1;
        c_cnt_bypass_en14: string  := "false";
        c_cnt_in_src14  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en14: string  := "false";
        c_cnt_prst14    : integer := 1;
        c_cnt_ph_mux_prst14: integer := 0;
        c_cnt_hi_div15  : integer := 1;
        c_cnt_lo_div15  : integer := 1;
        c_cnt_bypass_en15: string  := "false";
        c_cnt_in_src15  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en15: string  := "false";
        c_cnt_prst15    : integer := 1;
        c_cnt_ph_mux_prst15: integer := 0;
        c_cnt_hi_div16  : integer := 1;
        c_cnt_lo_div16  : integer := 1;
        c_cnt_bypass_en16: string  := "false";
        c_cnt_in_src16  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en16: string  := "false";
        c_cnt_prst16    : integer := 1;
        c_cnt_ph_mux_prst16: integer := 0;
        c_cnt_hi_div17  : integer := 1;
        c_cnt_lo_div17  : integer := 1;
        c_cnt_bypass_en17: string  := "false";
        c_cnt_in_src17  : string  := "ph_mux_clk";
        c_cnt_odd_div_duty_en17: string  := "false";
        c_cnt_prst17    : integer := 1;
        c_cnt_ph_mux_prst17: integer := 0;
        pll_vco_div     : integer := 1;
        pll_slf_rst     : string  := "false";
        pll_bw_sel      : string  := "low";
        pll_output_clk_frequency: string  := "0 MHz";
        pll_cp_current  : integer := 0;
        pll_bwctrl      : integer := 0;
        pll_fractional_division: integer := 1;
        pll_fractional_cout: integer := 24;
        pll_dsm_out_sel : string  := "1st_order";
        mimic_fbclk_type: string  := "gclk";
        pll_fbclk_mux_1 : string  := "glb";
        pll_fbclk_mux_2 : string  := "fb_1";
        pll_m_cnt_in_src: string  := "ph_mux_clk";
        pll_vcoph_div   : integer := 1;
        refclk1_frequency: string  := "0 MHz";
        pll_clkin_0_src : string  := "clk_0";
        pll_clkin_1_src : string  := "clk_0";
        pll_clk_loss_sw_en: string  := "false";
        pll_auto_clk_sw_en: string  := "false";
        pll_manu_clk_sw_en: string  := "false";
        pll_clk_sw_dly  : integer := 0;
        pll_extclk_0_cnt_src: string  := "pll_extclk_cnt_src_vss";
        pll_extclk_1_cnt_src: string  := "pll_extclk_cnt_src_vss"
    );
    port(
        refclk          : in     vl_logic;
        refclk1         : in     vl_logic;
        fbclk           : in     vl_logic;
        rst             : in     vl_logic;
        phase_en        : in     vl_logic;
        updn            : in     vl_logic;
        num_phase_shifts: in     vl_logic_vector(2 downto 0);
        scanclk         : in     vl_logic;
        cntsel          : in     vl_logic_vector(4 downto 0);
        reconfig_to_pll : in     vl_logic_vector(63 downto 0);
        extswitch       : in     vl_logic;
        adjpllin        : in     vl_logic;
        cclk            : in     vl_logic;
        outclk          : out    vl_logic_vector;
        fboutclk        : out    vl_logic;
        locked          : out    vl_logic;
        phase_done      : out    vl_logic;
        reconfig_from_pll: out    vl_logic_vector(63 downto 0);
        activeclk       : out    vl_logic;
        clkbad          : out    vl_logic_vector(1 downto 0);
        phout           : out    vl_logic_vector(7 downto 0);
        lvds_clk        : out    vl_logic_vector(1 downto 0);
        loaden          : out    vl_logic_vector(1 downto 0);
        extclk_out      : out    vl_logic_vector(1 downto 0);
        cascade_out     : out    vl_logic_vector;
        zdbfbclk        : inout  vl_logic
    );
end altera_pll;
