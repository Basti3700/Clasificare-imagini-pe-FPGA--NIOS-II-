`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BDc8F2taUbralhMgOjhCWU8ylNZ8hIGcYOjkpGdCOeuIwOttslXr8fr52lKocTH2
XA9nvmFhU07pY/f4SafAcAHWYSpIh/M1rArw2W4Apnvlat2dl60NY7nKf3mwOXf8
kyDwrflOcL311bu1x1EttweZqOFqvayff1RGpHpq1+tLC03BikG44tQ2KVEk/HTx
rAqMhNHkGEz1ka6HeXsp2SUuxdBcbddbW7pZkeSKStAjndaxJVG+8lY9+aeX8AvW
`protect END_PROTECTED
