`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1oNui5npD/KbrICWc2U71BWxhYJ5Sl6h5iHKUag8+0CrBOQkNYGK6CZwTwFoVw1
CX3lhb54GBodocBoYH+F9telz1qyDZ0VwiYcYF2aRgcl8RgL8dGO+jAPfTnQB8Uq
TMV5W/2nvjEtNABOKKI4/GYcQ6CkBGsy7idS9jA5BBaUbd317qTF9qzMX6E588yH
/uIbRIr1Mwx2qtZykIL0ldpQwEY3NN1gdvxl7q0ymYgJKh6X5UaM7J5lJdxCaKSs
h/7qi47GTNP3nOudotf7++O+gWNNlm2vhTu8DaJAcwG9M4WnLzopxkF+wn5ye3BJ
nalFTO8KtyEMmawwFWg3XmfJ36YngcWURtwSeUXtFsgCyLRtOGrJ52moz90MJogB
DcKafVWT2EC8BN1tTUSw6kvFKNFfXW1ICmVB4q6D0NYmQk3HjSO+7cPz5wAG1RTm
u8h3UGAJgYH1WEAO0CXrn5rEhynY+8w1BBOuk+L4tLeJqehhXS7LURcP3TIXl0u/
o5jXgtX0iBPfc1t1gzWnH2dKo0UzQN/6RbY+XTCT1q8sJzx4DIpStD9YMq3t3Wzd
8fOxBN3niB8wsMlU7pjQd0peYxiwISKWS5UEUGGEMfpJlrdrHL6Bbd/N8mQ6F8M9
Jc0kAalQXTHq1SkPHapal8zvljIcFRw+oHBknBrzG1h1+kT0Xrkfryy5ZqTm2IWE
Buqb4VQqoGAfuwPLqO1+Ssx1VTMh0eQYosnAvH5SRcPkHIFD64mSUNjgHrn7GxKa
oLa7RRiIpPzqMWmuLB6+mnp3hMGx0BbY5PAqr/QzO+0n1ri0SwENudcH5XKKPxFk
yvnCgTM7gMy1JcgGDfDKKtQ+tivrKNn7iKwd9PjQJVMO8/+7QjajJ7hOP2BMWmRZ
qjOXRkU4H2i6R/PLO586l2li64XqLg9z0/d48w2aDIEpGi/4TAE1mRU5PAXYibnG
Dp0QWMraEjKnLCsvaZbUGSyf7IvkfkT86hM7ayfCJObfNMqXJt1B72DLxklL8TTu
nMpYmZb6muwKOW1aT2wTQj3b5wNU0hEQCb0uJFvuElu4+WOd5Up6zZs5QZnbMvti
h9UAZUHi7L3nswyLfWz6FX1UqUW4Z8bTxyNeP+2nh9kaO80Dt59veWiVrM86684D
/DIeC9rIwIBCkkCXjfvZy4VzqQWtcphVLy4pgMBlQTIfUcVXT8OkJUZ2CtHjjLB1
yHbnyqNJ6ZG2xW07TbL8xhiv9vQMEaZGW3U/j9CHPZ5e4mqej4PRrpHVi6jUmowm
fAlVHd9r6fzdSckxqXHoncUQXpSSInwg9SvGPcOfF7m+5kQ7Mvwt4qZhZX5jjNKQ
lIpHoJtXzGtDL3ynFk2lMPo1GEcL+RQcgqlfQUOYpD7Fuo6TW08pGOrdwe8EZ7pc
vA4uUXQmJzwRHFiVnCyJbw/yGce0WCvjoNHgFODHULq8NOfQ/faz/R0GPtbyhAg0
8YvTYnFbFx4ZecM9jmtrZk47l/hy3/Fj8aO0B42Oes9JHYYTqjfGQPYxQQ5kFDh2
6jKLJEp0eOzdL+7yImKOJ8psiLT/2N1PED0A3efuzfQAA6v6l3p//BMIkUqeUSfu
wf4Zfm6snihujgcxXTOyeE+BlCKYpPzUN7YIemDXUwa0kWfnwoFGJfJZdrHHeAt0
6cAR6Val29OlhgzahHBbOvPIk6Z18C5UAASQRj6IHFa+Wp/A5Gs3dBlRGgCS6KvU
QZDzkH8w49QcoXn/zPEhzmz3mxPdrhbLV59Go/y1fhQv/X7eAENxmXJuCEncGgl2
T0z2PzLP3pUPutsaUQC4IL5JezMYOon4JpOGrdxh5ioO/XBjbe764yo3QMwHrsPs
KmQ/3DVkcUjkdVOcx17e++e0IRSxAgspTPbQCm//gVHoTJkQvfxT1/a+5KWLWtFY
K8iBy3IOhHAkTc+TSItY2r7qM48P+QeFnhR94cyl3zRsEPppIkG5WxaLfbf5MERl
gtoprpsilOQr9qa/uCuGzl5OL7PPtxuej8AvfaIVxCxsEAXnu1h7tn8TT6xIuucR
k0etrajwgLnVi8FRfjPhug8p9KWv3yKDAXI2XJh6DweVr0e2UOcn91m07UedM/Ta
sO+ZAUq6MKA31fq2UllIjvuWn9qQnh0OV+uYw/n9RtoDAB19qN+UER0I5QiH90H2
2Iipt+cv8KfdtyZ/wxvL3KZmGC0JGUJJmvWfbUHdtRQOu5UnmcD2QHCP+29heIQH
ri6JDu6T4nvQ7GbdyiOyCKZ4HLyHSMjCaoMjey63SYLyeGZGwn5XnQxByVX7uFcl
0awCMk0/ibOGVVw6ZWQUBU2JVcyUM8sFt20s3qkS2rhu37qgY1ThG3S6gtVlfp1H
gRbbhoV0xnbjkwmdndUhk3fPVBK5IsQrQ/NgvZuLnGiJThYwAzODYmMefSr87Zqg
iJuufujem113oDsgv6o3tubjuKuMWhVST2XhhxYMbPc0GHB5DANp2v8JKGNHDD9Q
KNVsn6vMUXcA33EHtxg7u/6UW9yxsiiM+vPU3qsjuGbUzI50UNVi0HTrpfPWkqTf
2GYpoMesbO74Eg+NLzUAImXixzDetSeJ//X2Cd9YwXC2kgNI033U2cqlzDF8N4MK
TUpK3a6t1DYQqVz7fqaZB4fUMp/UamMcYIoE+7Xm27joXHFwhj1TWnhl6UIzqCWz
QVrHL54RxQFzILYoDgruczMCb2aDohqMmD22JOQZsKZ/X5O+j+4vZlpFzqhhsFGL
EaWEhnnb7A/36aijnL/uezsx/Kv3Oj7sh0UyQr6KqvcehygaEC0VH4t86t4QKWJ5
s4PS9b+wcKLncCNE77AJY1xD8waO9ggxaKtNqJQQq16Z4qPXoUE6mn7qmz8lM4ZS
Bkqq5eM6VkWtzm6c3SX7fb8LawENP/Q+UeC93q3RpxcO4eDsDpj2YQN62Zs4TY6Y
7/XJd0p5AijyXt0rQMpz79sMHFmO9GY+UF5zWq79S0WnAQ1phWwFku8n/GXUzeEz
kzBrhCZ5dd3dWxrvR5BUmkMt4er08HXG4oim/iSjKAdZ5VuLMxIF3XtWt6y6/Ai6
iRhrKSk/JrLPmdE3YySOGOpesUGPU+RoYksJcKZ/HyqPaFPZm/m4yonWMQeXjVMz
32lXFbFUhkOjAQBGZiPPUlrVvbB1+fYnMuHC7fPAIqj/okCnmQqvPCr6NU/Tr5ro
CYY5pN6T4fbVgOMl+DTENvyPX70H63moX8udMeptfAnIeB4HOwyTqSckJnaONwlo
aFHKciPUzwVjkr8W07yhj6Gf7E/izODvyba39/r34JtmDCIEekoEozWYcQ8sf7Hh
I/UjlzkwI5AvWZ4eq1Ck0xu2Zxlool9oOfDSjC7aE70ZWGCkIU+lr/l/F6ppuC6f
Mr8kkT/mlFtSFeP+eMfgSVvQRiEGtvowAihwNFnXxSNLOkLstfDHi02cPLdbD+jL
G9N7750p/bXZTnXgnA+YMl9JZMVFc7q4IZ+k4bWrHGXwIXqzP/AAmLOQU71Dc9zl
0SntLPy2z+2JWz/pFU6HWJ75308twibP4jMao/9m6vZF6eJHy9bzscsis5UO/BAo
cW1oDVfdcfP5c/e9Kz7QY9cZ3HLJeU1y5HTkX8BBozwoN65eYXihe2I+iPQuTlob
Y/BoLMUqN/ItTATjvlj1fyOtlc0NTrdvTVHn5l9OopjWsen0mR48nNYRiRHqYP7M
CgOe3T6D27wg1a5DUb2bm1G+10Xn5QMtmXhgQwSdS26FAFh+VRAfLwqvdig932hX
zEN8D+VAM3M/g76KyIVKPIZ5JXDT7Ge/KEPY0XxUmq+0sc14rhnVR1rVVldtVf3W
GacKb3qaC1VRhbRBPLFdsFcYZ6To0axfE0iqclY7CFHx1LIIZ7o3y2wX82z0nTYY
4KV8Qp02hH7WoyTWglHhh+q1rZpSdNhgSXpG8h20JWKLeG5uWHVUL+ySKWV6vz9E
NnUkH34n/Md/bNskApsokEMNSxgeHNXcdhTL2m73bka7n2Q6oudg91S2IOsUIlYL
OSglb8G4wIzX0UNcsbvF11+E1e0tr5oHwLKMERU4pHmbSODK5LTflYL4LFCuuYak
KTe4McWeVagk+SNlm01CfhFn/rNsUhHuMgam2LESOux4MN9juQnOuox1DDQWljye
tUUGp7pWTyntS1ubboojLYKlzZLmBECbUDMvNAaFrpRU/RQk3RyHEX8i3AyjZhCZ
Zg/6pNwsC98QbzlP8j5Bo3bINRy13Om5H81czD2Gg6mHnyKjrkfnpUVvxj6Z92/t
acZubJi+ez6FDhgrPtdkw5Dh7+JON76EjstXM5/fv+0jJO104q6kv6t+DJQWMd5q
ylokYSdpORjzWfWCKD3SFDxEXVtjggzme++WVY8ttskQ5GLuuZM0/mcb4USkjtoZ
oVTVp5ezCwPb8tIwaoUQO7Rz7ChtrGAVapYvdne9WtKsRwVhPjJizWOPC5F3boCU
fTp9ehav2knVIvzibEVkKNKmi37ilsebyKgftNAa9NBHUJ9NPmSNJ49eWwwS3alx
QZcSeh/m2R5PbRZllz6uKzLdPAjtGZZse22NLoYyuyMhDDd2cVvywImjne8XKD0t
i15ggIPNDgQjAXzo39lxXFbOXPaRaaOOBrtukMlS8/u6PeptqJnUz5Ssx+z/bG6m
1QM4CbGf1kN/ZfbSpSmG0dqLU0uKDwScxbKE/opLtqxLr8VNRlNFbCPr8Qg/uSFU
z+HZ3UKe00qnxh9oO6X/a36+50vC1I7FbqjsJ2VAMAbg/coFJhnPqlyJP11fU/dj
KvUl0UFFlyJHxhtjgBOHWhkY+HT32nfzfVmwRaxNyH23OV0O/tBdBMuCfs4rdWAp
0yG385dpLI8NcBZR2TKH7cdDMoP5uSk0kTeNB58DRh2Y3tKqYIuPQNicqQNaB8NW
cKrN8jDHNA8khgKQT+6gypT0uQr5cXe8N+HYsK3P90rI1db/T90LtU2Dz3+vUrQl
MmqwISBS7R8jR2n3l3RpwVk9ViF/66HdpAWn6HtyrckS1db3vsmGe+bj97FdPcjT
AwluJRBQfsspN1tUguXdNhtWy7j8h/ouiXcYby736+6akTyCLSrof+brknRAFwVH
zH9CjOoj86Txao3EvSyq/vSw/LefZjPUQgWF/38R4qSlrKDZNePKY1KFpexOVygO
o74ZZyzYpMByxjr+pHJbPVJ4tvO95ecTktFQftyNV86hDAFqZzcTXMNuXgbdJ+G4
GtbI4uJxXsCNFAoSDlvcbNeUFvey04WawGYti0IXvOuC0rE+l/46VmGl2hUtBQZ5
54MruoAiuIsaSB+Sl9EmioCLpAhnQ64RXBeZV/EwQszPcONuoRYJgWoc+ba90hl9
2FHEoCRFh+h+ouJybuWs2twuP+TrQ1YaVXiEN9o1I3IeC8IfrkUk0Yv294KG8eKg
yA9Fl+rHQvxS0KpB+WRhtgINgXFZ08eMy04JrHmuI39mbdHeNJzeZK+Bf9YNCbWI
kIJdOu/emhWZGxCw0UThfLB7l7clS/Fnr3qDF3yD7a9YNMg7xYx9Zx0/b6URtudQ
UzP3jrzudBEEH+5n4ESn/DH2JTx0tgdGytfCoqStK9b8xBHS7ZyBkFnkVkpYxEo+
kN9UdZ0HycpSumswwHQI/ywoJ7AJyaKKTdZUvDAiEN9so5NfW2P9joXmneChFvlb
7ocb5K9LCDh0kl4vhBQihhc0B72Zm9I4LcuW4jPGypgZM1hp2wAZgMDBOWK3ESDW
HSi+MX6Ez/foOM3pTMZXQzjB76tcgp70UyRfKdgM275aehoyqXQJhbkaa5CTvvXY
KlKm2iKIh0yCcc8oB77HDjCz29dIHJ0lJ0dA/cHBiPcGC+BnyWuUYwLiQQy4+5y5
XmhxsNDs+oPWy/qxiHXW607yZHTEa11lwfzU9bLMK3CnftePs41AgsZQdKAShuQs
gtIINskac/BStqxsHABoyv8CGrGY9m6TXfNyYOQxR0pkGChEbzRqkbmzzIHPmz/o
9QwWQbUQ7hoTenf3Gbw5X8dt4vD2N4rMOfzjD+J20olNjTa9MqBuQqFePE0+eiSc
Ft7Dl63XiuytUQs5+X4NGP6scBNDlsVazcKd/m83eVo0hH2ZldOfhVl+aFYHy3cV
9IIOEp9IX4tb/n6pOtDYeFMrSJJ+YN4qcL0o0fOTduG8U1q5545PHoajnGvlJpiP
0ijOH/3o6WilmeW8+oYrf9bNODVBgUS3HskZdYWFNxC79ClIx6Key7ca9odDoK90
gDwBRrtD/OYHOV7Iz61tfg5y0aI+QEw63gYPlIIAM/Gl5oSp1yfEhT5m1Di64Yn5
F4Va54dJ/F7DsPIMNFICMnmlyG/3V79FApOi/ecS9TBpBzRGRgtnDvQKZeMcyIYn
x1w/1pemfOiTKOcbjtYpfWW3LvP7V0LRH/Esb8TLW8JQq795EFvTbePTqliSgUI9
gX8JDsLUfaSNNOiMaBDsFt/WnKfwjFeqZkjZmKAgHgKA+wBCcb238PVnJYMVuFzO
UC4KIZ8vnVvlquvkRJHT5cIAKtG4rRVM81vYuMFRleSxXsqHlByeGWVjevxrOTwK
oKvHBoG54P/rf+hRDo4+Jx6vui4GEK7TlBL0HQ7efulvddqdbA4FbR6FJ5XpsBYa
ATQDERHC73omSBbU0gPe8KH7++xbsPSPWpmiEabQmtPtCNpBXLnNBCN53+Lp0kgM
6xQEe7mQCJL20VnLWzL/btlScEfvlxGLTJ2ZlHvhRsRCt72n8/74pOCn0ZmU/2yx
TT0Sf8UhAMeAbFym/QWC5g==
`protect END_PROTECTED
