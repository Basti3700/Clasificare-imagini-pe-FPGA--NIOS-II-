`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDzf9CSn6KF/dSGrDHkY/m+q+VjRT4nV3F2CctQYpDVHV9a0+Zrsb0RAZwVvd6PU
mUAo9Ueb6jL2bXls2dm6A0p4f8UBDE4k8KmNQ9uuJNTga2vIs4a3fUG9/HrGZwrc
5j06MT7j8N3Vu1e2MP4FOE/HRNFFl0pWAGfdcZqFZGg+Jcz8UyvIzJyX7Kpl8mh9
ImdLALqLswhgGiwR7oeYulyHzbXqhTFKOGEngLhb9Q+BtAHpBlb45TNTgA+HvanW
pY4ke0YJ9k2lIXhA+ajCKcFaN8jXXuseHJFSjxNlR2adORkcvAR9nxyRwcAB7Zkb
tFmVzW+SwvVXL5FyPUxiwHpbg1/+Bgm1naZWkYJ+CVo=
`protect END_PROTECTED
