`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLd67EwuXgzMfuPhZGsVBlNvQ+VskIb5E30ZjuD/7WD+WUTGXiy0L2Ulz8Yw/Sx4
ZCMv/7lMgsw19mdcMgODpmhbAk+zfqkOKE9qT2o9Z1ba6L2VrQKR0tB96EBEfdla
LuiYV+1JbB9Pf3wxamIsdlPnwFQFmVjuls9RibbBYCVZa9TyuSgHLSWqdOv2k2z9
Qlceu7J4A8mD9QCfCjr2/kQsjZtbamh/nnFlsahW9JB+GZBpREZ3O1I2PaKQSVHa
oGIy9WNy9X/nNrpCdOrJ1J873M53lKtM2OBsXRPPvcq/8mrFqKWsn0eKXU+44Nop
8c9lOnIjaxAIM1WqGZILl8QFFJCT8/89phavPXlQrU8orY3LT7+nyULLdBkVHc93
`protect END_PROTECTED
