`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DVfDqO2Hdpn2vfvwERxPeRDGmHx1Fsz1Gdbv2SVfDJC8EaWY6jD4Wq9xjZrNy9qz
ahW7hBMpZfA6x2GRoOvhWDOl/8rnD432YFOVQrMhJNCni6i0h3gNgSIrKpsqgSXv
9t/v9Q0BBmsKR5CaNepqEWe6viRvoXU3mJsoG88XPpCZZ1IvGQeuxWT9K7SHa01V
adsvyG4oQjnvRqEy3sKd+cEz/ps6QcCEGE6cCEdmrp+aJ9/QxAJzoNOprjcTIbbv
M3jjjb1GUSl4M/YQvPbfS3kMa3qjzhQgAKRlHrr+ggrsnB523cxRBArSnt1i29Fm
devvwkNKyIACBzLZ9lT7lXjIRwAt5BjsU7wvO4gMBri2yNUb4bt+AIJLpA/AatEj
s8wdQvVIb+PD6762VxkbszWkRiLeUY9VAa9QEc/Qccz44G4A2/h3YFD2NE8dCCZ8
j5k+tLufOxuaVxinJJdNOgeNuPlZAWTMMGZ9vBF2PIdhnIsGGTGj9VBaV3c+Crs9
LYudXcdElZTkkRSeJbEi/WH2MbYbawuOYS8nlyYCSmQa9VK9rEeQwpSxukGf1yiC
+P2L2TTuVtKhfT8VGonQWlqIphGnhuq5lBgvEi040d9KTu7nozw38tptPaR2egxQ
GI5HRXVGGqX/X1bIQ88Ca4UPpyp144tNpJTbRlghSrnKHiXAU/DCNssxHaarRiDX
P6KaQGk2xvI0dN0EGsblI6mwqHlnFTuR85H66/DfzS7eVbwFtfXwg6misPszUQs0
aDjMb38KUlnAvXki2kXKo5ewm2rWSkqhJwDFmk5Vx8cZWt6MW47ORFBIJ8yfxC/j
QJMH/M+EqD7EaX50ZmstgLnPT/V1YeqfeRohNJbY0LVS06kC+tGiPF9E8QiOmlYw
cB6uYbJnL6WN/5KhTbF8am+KI+w8CWzDCwJsYn67viWI74VFVswPsTE60xbFZgyh
rHLx8/+3aPo1fhIGsBmLjGV/9Ltqo0kF2stKfESBx91UyU2PoJb0ngF1/fKACvtr
mtFFuJTOzahu6S+LU+DeocMJ0teru6tcFizxHbI7k3O4aUWV5eXLnHZcWTiNAluE
KQZYzTTVPcoBH1DymxN17KvIwY/xvibQKzIdbuFQPcY/b1Q0BnZX1EQCy6K0IbTg
76A9WYrYPzl42w1DCv7bjp9jJUpSNZYfXdQE2k6MiSFD8aLz3iqcyHI0vo45lvKI
/hy0YV4ToeSldZfMTlDpcmw4mcLTwDiMF6K43mDtEZG64i6qntM0n57a9kj0n2lo
OrAtd4t+t6qa2sLPc9Hc8ng9Eaj+gu9lpg9TnHTJgvPj7OUCs52kd0XiT5lN4vnr
tKiP62qwwjkLjUKHvpyhoZlRM7ObJlKD4ssKp+0qjsbJZ3Q1wVgxAneicVnuMnWO
f10rzhufqu0rVh/MvHq8kHO7sw8ja5kPiGhK7gjyQcQGGr5RCeumThIJpFO5TcNR
Ye0O81J/SnfqIQ0xQWwB4iucIN6G+AUdDPvbQf6MUN5YLtEGU9O0NOnrt/DaycCw
+g5NNFWxbijglf7uq13QTnQxo5bJDWLVN6OOcxnP/iGstqwqLXTxmpQ2/2vHvuUo
CHpOAe9gJtaePas+sYGFEAeZcbDbuk7DxFJ3VcFNbGr0/vr9AHrm6VGOr44pQB/E
awU/QGeKvKpXhxS4ECYn+uBp6Tp1U/c06+Lr14TCjcK4DmqWk8BgfWe99iRlFS0C
cUsnXJF9vGit9O4M2W4o4u6nz/kPj9Rb4eZSzy4kY8jF4A6SgyMsTC0WX+y7gNaf
NIK1FfevLOVPHsvalVq/4ler4EyPtJVPyHFWBML7C18S6TQD/GmL3heVZgAum9pw
yfgmU/53eoV49P9beMj0JMohY+eHiEt/jmB4Bul7sTtACYSEPHYH14ReZdXgCP/L
VYYcBfbOoKABTkGcpwsgCA5A0vt5fSsLrzzcTltkFBwqJQxoUe543dwzVj+j7tsp
drTQrtlrM45U9Jg3rwvz9qDrVq7NhtasPSjCj1cE8GiQiTVVmi7gjEOcRwqclsmm
LhxjhAfmsZQsWjDYpgSm/icvMsnL5YADtDq6um8vxEAEQqlUQrDJ5ynJoDSgQk6N
q2ZKgxY3mmRaNh31YoxGoZJE5g5V1oq0XrYyQDnoVw2KMv0se2pz6BuJ8PevYovz
KuRuo2ZJleeswBofmqzAchqgKhD/Q8ThHzmcDLWEMPs+hq0/TSvR1PyWO2GybBZ8
OOKAqL4NcV2f8MYCTI8qUsRNNr8MorpjUe3QWrKwSa37mRrvbIC5C2BpcTSN0y1w
l62soePjFu1L1oQgaXpe/sApUQHhQ+AyHw/ML5U6IAXC+NT5ywnm9Usja8Wyt5Me
x2urqyUr3M1AGpwZDjNurIwJM5gPGcZqyejrWpIkFf2jV4j1ad/323+qOn/D90r0
0p8/GTqD45U1IDRbhQsqyv3pYfXyXwjH9x0iRRPDodDGiKh6ODuagmbPVqhikmd/
Zod3lq9+3xNcetLwp4pqjkcELaT0uUuyHjPWC2EWCFNhWSzkF9V1q7dQcdUnok7b
ssVqD3nqi3OEkGte5FoRRq8u2y6yhmjuoKTSHadsqivY+T+OBX290O+6vKtmexYc
v6sQxgUYxRi7nZrL9dTPWSSXpkEqBokD2DVhE/Q2Qmdi3iZo5d9zX1zb97MtM7fD
QFtRRVOr6NaCIFszNHw/Wa7HsKMlYx/BxC8N4geiQDmr2ULioYGE0dJCPrF3wDvO
E+GYCwEUyyRn2m3FyExlRkjZK1309tS0j4VsWrXiAHlxPtEpP01/r8LPWudfss3V
UsMW6YclQoy7NiBd9Ge9GVamc9myBSopd1NFklvhq7gm+chRHtAutqNuQl1Ygh9S
rwIXothn1PtOUI1CRxxWnwMjW4hxPgR6tbaFYCIdWPL755+rd5vm1wTIebDVemyL
aUu7QJcSiubvNZ36qXBTd2MdGaEVzxgHBfwBnkne8aMPmyzYQ+4kFPmdr6QCWi+T
gHvvc/7wjAgbJYMMDsqdOk8/BEKeEGHp/V+1HdP3QqYqY23DI+M/WluPjxi2IfK1
uq1yHOklBrMQK/TMmmx5ua7LXPSI3R0GreYWhLb4x6d6QtbgqCP+7qQ377iRRubz
VNyXhf394w8PMDGlZJXs41YrA3fbF6zMvlvyvmnrat/xS/5r9thNauMQEOfMm1z4
0NGmQk+Rw09gzk7Wgf/JbOP0JrWS5PloY3F9il1iJNbTTQKLFRw/3QPHJ/Wfuq20
KJz+KCaX0d/+Wsf9PaPdSWXZeYlYmCp2E0l2pvfwWu5kD3BHFsmEhzt0AA8+NDNB
BKLMnvDtxjTxIyzSVE3LWnvjEBLIBSwcWZJvMq31OISSTHM56xb5xY81OIMVB1Al
n0GbqgltuW7y4vzIyXANpgeKoFfqHWnedTV54CfNh031aA/XcxJdixkFIlhVV+BR
Lp11F98a93ezQ9xvQ0gAbIDhTg9D6G4HDp6IlphHJiIufUIWaj6bsiLafAHqjCTT
+8GIRRDWQRS5Gpr3LPKmBd9zKYPrvytsh2HsWu2KIefTVCeMnzo8wDK8yL7JBXpu
RK4Ika+vxvQF8YQgYlTip0ShfDVQWebslAkl//lBo+rbI57xeNpqscztpq6ZBGn6
oLToG067As4U72uPPmlTcbLooQU/1jm/uqXFas+LI3TZQXT1lpbIXwOIAYuKR3GQ
RDXu7/TSDDvM+40VA8kWH/UFvEy1zbQZCdQZGoKMn53SCoRBEuym5zRRx5FFHrmQ
LxKYbvX/BtjYHmiqybLdCM4nqgbhW4EHZ5dXVTXPrMNT8cC3OwwppavsX4PaNXRx
b1mPiEP13tpfNTK5MZ7BM0UA5haPG/nkylZdvM5JKmNwRQiaISKKbS1a3tdKQzSU
FyR5K0UBRV+hAtji6SJnXyBGuH2sAhgF5/Cpq6pvbRXTK9YYO2R/IvqrQ9JIPPpP
/DS/xooEcCv3L33OGByhEpT8QmB61QwlKcCiWRX3KQwAR0ws77tJiNpEVYcfc47p
VaqF0JJc67uBhv9u2yOvLq58rFtYmARnVRuDLyMJx4iIlb7Dw/O5/5ILOukF/Yk0
g45OZqR1Dr2eVHbVj2zSKwXmnWtoLMV/qdiQ0+c41oG06B2byGZ8QMKR+WX1I2BJ
aAocnSUEvKN48qwc5NoOawIoGHur706FEXomA1/RUcKv2+nHb0/yEs0RDzOUnVw8
yVjAbn+MpPmSaTXU3BvOnlAfZ6ZxCN0/D0Mj58LnN+F1QhC6QFN0UrDG11dkIltG
rCLyPB+9BbsEsn7nyE6pDtOPNrfgHLEnAXFu7F99Vh1klTJaD2M6FoQYmBooOCxF
elDx9lFW2q4HIEoArME5rRTU84gudEFVfiDWJk5C9Lm8X5Zns5byAQgjonO75Ti/
`protect END_PROTECTED
