`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9/GhvclvUhdjvZ96b/cOkQpSBdFj/Br7VsvXgElQaTMBvGYh6+ckMRL9phHKpbx
xz3X5SCo2N0ueE4cEJl4rCJ7VFOZvn04ZmngoFUCWI/ou6R1J+QGvnksMKpiyA1x
vF2APobZVqKOSSVYFw9lD3mqRYIgCb8bc4jTLq7bu/FcGRf4qN0ZKoUlNdgOJJSI
RgodvK/tCkJo/pI4gZJdi8MLn37P1xPPdGOPD1TqiZRaWdnDc+0i9O5EcEvWRG1/
yG+BzQu+OdCxlS+Dzs1SZwhFx6U+8on83Bf1e0fum7i/P+Wt2jFvDps8FRGGjsrd
edfIsWsamC7vzACYHAIfSIuUjyjyVvloOTHsT4Z455RXwKAG4rlqiua8VKfcFW00
jh82oWvD+lJVfvnxCiiCskjIEuzv12c1G85Wj/khCXHj9sUrioh6i3m/ln8+OV24
KcZNsqKp6gwuV5lVVrZCocOCvQnU8XGiSivgntIh3LJx2bglgcsyZRQyENG0SqGB
Hf/+/7N1ao9dunpdYUDPbiCGoOEIm6ysg62yflJcKgW94owz8ZnvREtqMyrYywfA
JLPKuQmE5TXgV1ccq6o8jvpFHXbm7QLtUfWqMZkR2BBzSzRvv+2IQ/wCUsk7hoVQ
ooafqi9M5f2S/GJbAzEDaIHR3qS8QvkP5NBU72aqKNCWGTLWa986TpIhn3c9fqZO
19AC5NW41F+EWuT0YxelGe6yom57lt8TNtAwuXSaeqW1BW/es46IHm9OswClx+rq
EF+MHuSUpzEzsCEJ9AwJ2sv5NpteruWzb/UZVxkcJwrlMf16uje0jlEjQjLVy5gU
PjYNQN5kmnWl3nQDjAGOoH7gQBSVBC66bK0IUV1cbkpEoQZ5mBd0zBhL7CcawUE1
5juY2lb/NsfyxboW/lA0nKLtsUzqSe2wcoDUUhx77bFl8XvXKkNYhdh6WJnFiEcE
5IBRnWse9uaNW6qhPpRZ0N68aAeg0ylbdYHZWI1kgiDujx2o4Ovwfptwvp8Pj0Xd
FuhIvfDZG/dvakcw9MgLAeuI7pzt7dMoDAF4OEbWUXwjepJe85mtJMboYtnxqLHy
oRSbGzw1BV2TbvZVTmIuHE3HO32NrOP4jJLz8mg/U2FfCdFjJT7tF56nB9eznAA3
o9mGbFcL1I95zqKyq9VOWL9lPZKTbQcg2/arR+CB1cpVyD7umoHgJPoUaaeeSPCw
HAUz37iDjRPYsKaDWQgSKcEJrn9jAX2nZu0gzG5R1XtV7qRXaDvVYdYeWCStG9q9
GX1wrcTPA1SQ4B1qnIeO67+IXdMGiZWDIR9VxwYYihGNH0eGAHgIH86pdY3pz1bQ
2pd5ctVcVz2AiLfFs4nTP+9wNB+IOhFF7MP3j89wki0Y5tokTNdmeKrDrmWA2ZE3
tK0JjEfjkbQ1Oqx9g+zjLPhTrmQOPq2xsaYlRe1ksH8JxdNWARI+KwyLLxdRsb0m
FRDfHI89Y5ifYmyGCFRDr88jKi7Ll6L/JxyfvkDw5/Y2Fbhyi84KD6CMqn/NK8Qp
Ns9Z3MSVZFfE99lCgcgcnHpbHTppN8Ptxn3V3L8sZSnA+Etxc9nhA/OGuN8t0XTF
yGGJwfqyVgVZxmDRlWlg9mGlrpYOcXZ5MimBd0z6aJ5yy/VR3qqdLqVDk6EFkLmB
RQZ6hGX6YzkHzQjBoj3uYIVLAcBZniFA2SRsfEmEjw1SVV5aX9wl/zva3tR4pmsn
OFFkA4iFBw9iE0XEoHzaaheIAC+cybLFB2CBjAeO0yugoaDt3adnm83PRFqLUKai
p1Kle+iqt5/Z+SCZ8fBvTCElvCk5jZ86e0naOZh9ywz5uq6C4MWlYenrfCx+putf
IlvM+TV3wexrddIu6xpOW12vXa+dgNR/lVDGPDAfwjlpe1YTc3tWFuYyNO2XKY1L
q5/I0KzA52mpUDUjlRHpmMi2ex2GYVsKD6A5KP1cSBubDlcpNY4EnviqrfPXyAVc
5sKSMXWITIAM9p6RKne1r+wBXFo0iAWfJ9vNU5Tu0AqZWzS/lGOEAfPhLsVjqDbf
3ya81sdFD2VcnlAvD48aXU1o2Yee4DYhGwYERzh2bGB46I09t0t/imP+Z4mqZ+Z6
6BidmEFefnMlgNO8M9tn9Mw7HtEwyi3k9kiUm8SaUe4/wI1IRl6eyjN78ZpV3cBr
QfOSl65YUEvwQEEUd/6P7rSAYAN1bxMBUo7A50qxNFQGz/FR/W5ocjaV5jCbOJ60
g7HfcxOypKfmcW9fvPtqV2jfk7yWON35lKqXOVNuFv9Ddu6cZF2VEl56SXedCeTJ
FFL7TQRVDb+CazV3P9/K+CmWztBgS/cveifAoTWGmUbg82TaTloKG5vQeyaEy8S4
b8Mu1jVQT+ssHnfK438ACnfh8Luvs9wXAtpW5UwChPOYyf1C+YGVeICC/P/qByD8
o/+Ib3WQCW7G3D/MmAaFL0t7bQsZgFXRC/MOxdX1eaiVFgMP2IlT4nDSjX+ChDdm
Rf2kz8Hmszj3Z+Br5lRRdVTdeQYbRAKK6xcGXG4FagWaFA1l0YKVXqD3feP+HVj4
EfNX3Bx3rPqkqV5LKA4eBE4VGjti3YnBALUvUiFUKDU1G0n1tCLXU0W8ySBUlM+e
UjdXKSDsFyQmULwkRFVwgcFBXmdGLqi3ik5dmFuB1UfuvPhNOyINNX9pbOfbmEZJ
BLOv+jus+plnbT8MHxAVE/1RRb1aVG/VgVMdojkNmg08/ABrF97Qg1cXhxBuyUad
7f+RVHnp7SpC2FProSJR/rWFNr3xxeBPjqUDKrO0fGQ=
`protect END_PROTECTED
