library verilog;
use verilog.vl_types.all;
entity ama_systolic_adder_function is
    generic(
        width_data_in   : integer := 1;
        width_chainin   : integer := 1;
        width_data_out  : integer := 1;
        number_of_adder_input: integer := 1;
        systolic_delay1 : string  := "UNREGISTERED";
        systolic_aclr1  : string  := "NONE";
        systolic_delay3 : string  := "UNREGISTERED";
        systolic_aclr3  : string  := "NONE";
        systolic_sclr1  : string  := "NONE";
        systolic_sclr3  : string  := "NONE";
        adder1_direction: string  := "NONE";
        adder3_direction: string  := "NONE";
        port_addnsub1   : string  := "PORT_UNUSED";
        addnsub_multiplier_register1: string  := "CLOCK0";
        addnsub_multiplier_aclr1: string  := "ACLR3";
        port_addnsub3   : string  := "PORT_UNUSED";
        addnsub_multiplier_register3: string  := "CLOCK0";
        addnsub_multiplier_aclr3: string  := "ACLR3";
        addnsub_multiplier_sclr1: string  := "SCLR3";
        addnsub_multiplier_sclr3: string  := "SCLR3";
        use_subnadd     : string  := "NO";
        latency         : integer := 0;
        addnsub_multiplier_latency_clock1: string  := "UNREGISTERED";
        addnsub_multiplier_latency_aclr1: string  := "NONE";
        addnsub_multiplier_latency_clock3: string  := "UNREGISTERED";
        addnsub_multiplier_latency_aclr3: string  := "NONE";
        addnsub_multiplier_latency_sclr1: string  := "NONE";
        addnsub_multiplier_latency_sclr3: string  := "NONE"
    );
    port(
        data_in_0       : in     vl_logic_vector;
        data_in_1       : in     vl_logic_vector;
        data_in_2       : in     vl_logic_vector;
        data_in_3       : in     vl_logic_vector;
        chainin         : in     vl_logic_vector;
        clock           : in     vl_logic_vector(3 downto 0);
        aclr            : in     vl_logic_vector(3 downto 0);
        sclr            : in     vl_logic_vector(3 downto 0);
        ena             : in     vl_logic_vector(3 downto 0);
        data_out        : out    vl_logic_vector;
        addnsub1        : in     vl_logic;
        addnsub3        : in     vl_logic
    );
end ama_systolic_adder_function;
