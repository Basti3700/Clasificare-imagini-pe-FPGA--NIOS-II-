`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ykt56ty2GVTiCi5azWGLAIDPTQs2t8GeLk8xHbXq0uqC3cW2rcB4qPux3yoUypAz
+xJYlCsT7SMuf58aX3yQjAkTfQVUPqwEy+SBsiiEa1AEWcb8BYaegfYzXaxjHvgu
2xYyD+n/37z5I2Goi/l/OifxruWXfQ2CGpEhqaCcCJHQmKtF/oFEVafjrC1Me4AZ
tJuW+R3deouz3kzuMxzSs2qVrXquUSYkUc1i4NvLeIRbxOAL+AbywIfg35PlrXtn
1rwOguwyLXqZBHpQySSLmkydVEIodq2meTqv4q+uqaX6j6XPVr3gFG7LnQtcR0Wl
1j6M6pXIsKqJlib8nAAaENw2vFr2Kk5BLmzXRYNbUyqe9OiQUA2YkJp5fQOicYWE
WlQcMn2tofIfiSTrNYG0Pwt4AaWqhaidOZokwR9lAYRHzS4UWcTjTInIXMHmLF4p
j4vTwmVChXcOeRUYnvJqOTzDpoNPRdL6nruzbo+YOCtDwtM5wxICrqjriKIvxStf
frYfR+aP3XJAGnRecfG4DqaTcBPsxi6Ei8czxPqnwN4+l0DcXKa+If0X8kJNl/vy
8TQgVBmk3Leo75V8NoCycsmsssoAWrP3wLoOAbm89Mj9RsIA19qyNMsm/mOMvjYK
tHZGmlOWVF8j3B4dwsA6KowOp19aElQmhy3yN//Dwm5LDCJNlw3/UnucndT7KMLj
oS7d3+qrUuuluaH/Edk2uEKM3+jA7fT3QBw1pGtWPuNeeORcuJa9nf3r4/y2xQ+1
Pulc6ucI66YihwzP6XXmSjSE/m31bkpsgSjxOsVfOHH2nKdADO+IUv86CvEf8z7Y
LotUUUm79pFj+Qr9gIVmdOD8NGTtAWvTQGRMrGKm46L4u7n2TR0ufkTUQNx2HyPE
AhtMViCVrRG85f6SXzy1xvDthOOv/i/69MSo57QkCLNHCvGHOWx0N3zUXtuBFJlV
d1Bl/0YetgwRCV3bYt4TM7fa5RK04KQj6LC8DmOsKrxefVlcF/73Z42448aOlBcN
RaeP7MZ77dumA6NiC4aqi4h9SP3MOhn5EckxoIvWdyptaPhUgXz6tBJlhYB0iEXV
IGSnhr2y4ZneL5lGV2tbl1UqlRWdpv4W7POk4kgWHWykwVbhRhx48maZ7ZCQygm3
5I4rdWlihX3f0I8RTFTNNdyEsSXdaDh8TQ0LwDChcqQixFBFe42n1nLm7IpGp8o3
TJquYMebk84Wx8j0+d/o5T56XDxfeqIaRpTwZbS3i6qI6RPlFyCw2zJBXuuxQ9PA
y3UnGZ0SGVz/DHi9lE9FCEFySxgO/eEnHlt3MEDh9rWLqjf9XhusxhQ6JrjPFaZI
piHqWBgZiWyl1+IY/s6uWFis2t5gpAQZEMdX/xqWxcJIS4k4bfMB5DjeRRWI8bn3
wJcLVSqISb8Y/aWKmiHT8+XeVCkiNt2p4KthCKuVtE/OBVJ4g6x96l7KVZNOCoHv
vnhui4jlLAff1U+o7HbvkdJS71/zIZyLhOaWPDpIW3Ak7aHY5XYXVMJOlCPRu3RT
Q2GEq24RZrezZW5P6KQaufEmhYYaUY8WrHa4GY/0yRvOaXevZwUICOPZJ3Lnf5bh
fzZc4ySayE+Pq97BMUmCN61GF0BE6m93yizEMRfbTSbJugsEvHlkyK3dCKiR+LE1
sfXb3DUYGvwWoHzOz3FEcEnS8xoD2oRsvVED/38jajRGkIZ2QliQcKtKn7R0ZtI/
FLOIxQr+fulRBaiVVmoAErTlV0NrrxZyh5CqZ/Q0YYJcn1WfLEvr0B3MrzQwUNQx
TfksoKg/Xa8Jdn8th+9O7qG8ekBd+NKVbcR6/l7F57LyGuwAdQaygpDB0oZwXqdB
K8fPraNAsCsGC07NXRMavK44SF6IVZgaLD8wZ9HYi+4JdhXvSqnP1aUMXa3nWdsD
fdnGEniUD/S0xa6sI+uIZPAB+MbtyuZGzIVbtFZriV/Vr2BnF4B46sNSyv5jPaFQ
m2txSRCl91bshGymnmHaM0y5660RZpuaVTgiIgV/SyopxEhcRY3q/SVU+LKKcjbU
BuCHBcnXRQCoasGuNuGPhQ==
`protect END_PROTECTED
