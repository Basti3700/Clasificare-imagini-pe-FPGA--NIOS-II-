`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jw0BSBr1pAvhtMXFag2XzdzhsFg7fHLd2+lHyRm+SXOIsHuwLkdv3Qi7/XM8hcfT
wVskEa/QIJdsbli5ppAp3flQliwFrgCzdTQ5A1wLF/Hb8sbJ0qiujA2asEyubUdq
P6KsKwOWqc3vu9JdUrI/uoOoNAWhVordnaYbaiiz9SApEPrplo8uRHicrH7+expp
VDd0WmJ4ToZxPugsIubwufz+HvOGDUH9Pyl41l19CVPZ7Z+YoDl+aT8q/+ZJ85q2
MrGSSk3qu5ZwOl8v2zkbIqsaSmJhWy28WA0EEyJhr2JON+nqQ4g05v9UZfhL49QA
Pa8qKQ9+Jxce4RimbvQTb+BQV0tNXO2iXq3dX678Y/c5rSX2i3KdPa46b2wlvI3W
JUov2i7tV8gfmi4/LVoxccw4hLZH2Jh2zbZ6IWArDJ9LqaDT6iObSBmvrIJVU2TK
gXPY64jWnozTNvQbU7aJyxlgduE2e/J4selxuj4lJQ9ii3bE+qLhrhOYz8XtP8j5
CFfy2nZsJmPC7q90rF8zfQP4Qlsi0lYn2LvpauPz6TiHdJiQiJ5cpn+vlpa6oo/S
NzVa7Qtt/dx5tbM6aKnR8959HNPwskXvsP1j1onJZpaE/K2yvT2yi7Sjeduaj0Kk
FtXbfzT1vUFWozTgmpsIxEMNnYky2svaUMXGHp9yuMmRE0kluPAFQbtMk+Ypzgpz
8YBtZpp+jRDWmKlR2smUx+DyvGdrKjEYu2GPcfBGddIItZTx9RlcLh3JLKrnNRds
+rnN799+r+hfPdPaPnX1CkBPUNNdfNLOZpXvbxY8nW06VrZhjubWAuUS990uXlhS
HIezRp6+738mYsnbTujQE3yDRlspK51iQBr3liqyTyLDRZOKHVBipWjAPJPBpYK7
sz9NAysb5GWLgRAS6R6/g1UX+6mzYdCQdMab4I8/s08jOTR7AClE7KYdPOW44CGG
ZXMzxU0KFuqTKuxPzWUfzD2VYUfZArPXcBiezfnBhRtTZwmVOS/X+pjAOTya80L7
tXoIHV9VF1o+LjCd+c5/v8qaK8IpwyWbcL1jRQTZyfp292U0x86Z8B1AaZsJcr8S
/Td/e8s7/Xbs3PCtMnpGkWUGZ/dV5NCA8kxHgcprKgRHUjcmn0tk/Uq/VIINNeyG
jfxB9Lic5ijkjKVZydid4io/ET57E1h4BtvPk/rgvRf81KaBz9b48TeFJ0P43Pzt
tEH4ggsoOOPNnZ1pIeiEOayDNbhqE7lyzfO5rTYVZgfjdL1TBjOVHoPvz+uSUMTS
9dxv8bk7tlGmTPQ+GEDOPNZhQz7q0Du+S5V6phIgSOkO3RRKxzPV6VRw8sTiGtjW
KHnlkcu5nq6UZp5R/RWmX8vF889xtc0sCxU8kryAFuTQvs3YtoUTjvS9OauceQZc
LutJWXgWkKZcKlNlsOk2qYPE/bwRGIOugeuWKNAK7tQsf3MQ3HD4fNokzO7YC6uI
KaDhjp8JlWgsD+joZRoCEkuZcXf45WJYwAVRsLmObY97ne1d0aiNFm43KnpFdKM1
CEwpLbyPfH/rl6rm3rMLCx+wFzRe9HlHASGuAMRqgkZ6N01S+ZxLK3jHWnlWkY0k
An5zRqt2dKkzHx3V4pfD+8G6Sd89+1n0e1yOz0jPm4fNUz9lpYPxAOII7O9TDc7P
i4/+5hJTPj4GCCx5nkEn0ATv/EzPSiZGXFnOqSYON7CuMx86Z+FkczuMTFP5w4Zq
FCU/upaNGj7ILVlcBNPkCXKSak6NXGA43qaGHC2m4YiDZ60eKUXyMgQAAez/YPi6
sTMVu3ju1R9BMAgwfhGXknu6vZlSCqjIyZX+FuuSFEqi25bN0MkcS2F2ywMiNn8v
ziOzb4WQ4tq2OIPd045DlIqyPCxhlFzjAL0r0nO25aoM32OsGbOCg9LOmakezCy8
kfTwg8Joc+AkiHMfYKk1IQIoEIirIfwPCAXTkGX2lQF52+87oRxuCdv7ph5fTRGI
zX7mSpD0SzoY1Atk0bhyqV0IFcladWmO+IheoTo7H4i6HCLlV+5NqupsxobFKuYF
TV0j23/FHbvskf0q3z3l8NAUVZYIC+atZygt5AmH6D/38IT4UQ0+oMrg23Sx64hP
HVb3tYEz751rWVlEhQAttI4R8GZHfojw35VLeVaH5Z3iB7b5qqAJ5Gs5W8DExot/
J+c5oGT4t7MVjAIhCb10vL1kHhl/206h3P6MeELxNYjNMkpAF/mks3TUykYv5rf/
XFQHSSFWpZTVI/xJI8v9nWhMhkBb3W4G8SoF915z4nmZVBoYBjZ79GQOt6Ov2B7v
pr1Y/q5jEwakvAeOJfhnlGkSDudAyzuTaqAuiDwiF0DqKPIM9ei9aVzZ+WwSc5qP
OzQh1HG9aP9wQP0e1JCGqt4apZ8xk9ZxdS0qc1ImLZRbUl5jWsVIb3RkgDtmZX8v
UVDBKIebGYTQSYVGLtWp5iP5JYcJKm1dNVMvJkBbzNXGhLm+3/ud7nUPyozUFbSO
Q87xhi3nrN1gsJKKODa669rgJiVBz4wRY5osTzJX4aiRSryJcEKa9O+9Ys8cvf8s
YHT4GwRvwmxpPgINHusA0GYECuTfjbKkyDl+oCjacnYzqjJ6Ittyzc3bqDdiGOqO
a//lezQrEi8kAYgR8HrSFm8UK9ZElqeYJ2KuzYHA/Vrz4tr6aHit+bWJAKWc6+Zp
NxgJWvywCXZBRCF4ndwA/Yzv4PjgdihtTh7+8Ei5BX4zLExuqIlDDpp9dYJ5laqB
pTsZlbR8XVhNA0fo20q4/LbDSJZtyYfSMHWH1lMuKOROjpzLEO/1b0bxnd60R8kd
Ga5GPw9QiDDZrYk5vIfetpD9L2NR5p6UkuNh+Wn6Rwbm9OY6yL3J/cdv4bVZIuHf
1kvTHoYgYayk+JFRtpa7PV4ZHzpxWS8ZvbiCe/l9NjzobmMUBkQGiWhPl9VBh0dQ
sh/dY/SUP2KOkH1gGQlAuoMtohQc9se4cEYgPUJf5nTUXExuz+xLIAB4SXhwesx5
Or3pJJpLeiTZ9UQ43Hu/lcr4gA90tnVNrUnFqDpOe/M5RMpcBjewRrmmfu7G0qvw
gF4C40rHtL77cwSvJO12drqpEIpx6iNs2kdYZaykYK3hl6op2rK6S5lDso4HxxOn
Vu7d3qlB0j2KueBlHQTO1GQQkaMCBPpWYy6O2HKF88TQLTKzDMvgAHHDYhQ8CTaw
cTgjwtN4nd7OOVBAdG9FAtFbQvSw+EfgeAxXhJQizSMMv1EJMmY4rClsXL6OuHfY
Cos05XtSZcUOtfuus2CxW5Thlz7Mg2mGjr2MF/ze0Kex0+kdAIIqdtlxaHhAwMir
am+eV/q33B5g7pzDbm/fUZbdRf7xP7Qf2HbBh1DPcTUyMjyeAZ5Yo3csHBgK2Bh9
cSfToHpOEH5hPnMgdP/YyW+m02CLJAcZu+fVX1/pZ66rTO3sOftrZEMk+o7hwcJZ
RBF7rnx/FND9RFzhntE5APfn3aSwc3QosCIefe7tujRUvLsqcnEeOIzBqAXc6oC3
1lqoFIBVF3thfU7+QJvvrO4Vf1TOjmZGl/B/GFDSqKU1XZENE/S5PQ9T2esMzAfs
NPcIYpetOZc6NziW4RMthMgXRZGsCK45XbEMyJN5QJ0pXhGtYujNtC3frKfYm6zz
BwJCKdYw9XMmvwdeo0wdgtXjgBf6jvJeC/TvyWinUB1p2Upjv6Mmdw77OmNRTL8Z
1ZlD2TInpWDuG5K59zkMsiaVckNUfYt366RaSLwrA6VFFNGkF4i9cK8Wc8JmF1SV
i5C5mY5ivXazvz6+9dlAwB0HTSq7PuLuQYTWMnQJuFmCgyGLxPsFMqHNcbjyfbnZ
G6o2DE1ZBMDvEtVgdO7xNQzCc6XY+JrOIOloVllx3YpPpiEjzV6kTehIxPWbexYS
omu/tpMWZ3K6Uwdkjg0YZ6pXwWSGtcGTQmvRu+PQH+9YDaJ2fa7vR3oCbVfRWoIG
YxkebNju0V3b7EUc4S+6V64kuXEPmXOwfwJZG7DfJN4Lf7lP6StVaK/UdruwylPi
L81S9s1tDiekLBoMJlQI+hG7ldZs2rvgseu4S02Th3WnyX3Wt/lDZzjjBcXD5VBV
TyQMPA7+BcDohIeRlKQfdSn363mhv9beyq0HqiolD0rSgLhVOmt40QcajmTDAtYn
dt3RcY+TpUgsRcICyp5bEHyTEmOABE7W9A99MiTbDfbrzZ2z6AyBrLTqmBll9/pb
1Ds0yKMNmFc7KsNmwbnLb+xbycEfpjl251P1o/kXUkN6yCKxnQJwdxbuZwNZk56r
ar1zbUuyZmbt88Y/wL7HAap3S5iE4zb6MGX9qS7tMifJ54nsbjLj8BJ9Rrg7Ufu0
TApjEfxypaCpo7OVKjBmePrNTWagUtglnb7U3gxMXLMYUBACR4PG9hQA8qduDxnG
SPfWpwoLqGXfRLLBFKZaPKweXAxX8llri1ISAkbfsGsUO2nRRwQE9OQWsVfv+TFW
cVSxAuK+6N+OTs+/2S80a2pL60JHlFgQ8JfEgbtloIOmIs6m7aHLBwsZOwSwXqCN
/ecT0T0Jx98GskC4iMbW1Wh78eCAmHGM7v/Z71Gfb0ttGLSKgBx5DBucpOdcSBGc
bvWajFOaqz9Ovv/w5NKKbB66ZO/nx9CNEISIpnva/4gB9a9JZl5+i/ICm6XDiKYB
unKXX3elkLiJ1b0iwtOioC14LwWfKnITcdoI5Mu0+lltPBZ6w3fpR6+l4L3K5O7D
f62T/H73V/qnUIzq1jowdrC4yaGa0hSyvu5HR7zlgI7+JsPlBToqiCwxm8F4sCnM
SsAByKlBZQ7cxicutEt3LPbBwEthQ8vL+onPL0DaUcEhS1cOooYlOMa0U9wdkbpe
Mc44u9OwAgVJ05Wcb2+3turU5bE6dYJqjxqQOHiph7TGzjOYNDtaisvC7RlvF355
vIcLL37tgAyF5KqwC8uKcQB+xx8IBHTTv5PdThn3qWS5wFLiaF1V/DGTkWeKFBpR
bzkMpdgVW7Ww2DKsexCz0pH6C0F9PZPFvBr687JOMknNbFNItcJJyy+c2ybxzxWL
m/L/LBA3yWxYJzK+bQRw36pJKMIYaQbOworuZujyjXLuv9klWQY5o6N+Pq4yO/JP
KS1syADbO+aroYie9e4Muwzdo+AkSQE5M9l7uERIAHhIM6DrMeJK81yHH++KqrLa
I7VweY9R9VNherwNwNiMZoDuzTwlRWA7a1SIxc9KNCMpi7T/+HIP/KtOYZ4h65FH
Z9CTCLyJkgavucdszyojd7cT506Z2/DA176oL9qmVmdc3Joq8Wv+KDIStq2Qov/q
c+EremmpLTI5NgiZ7J89u4MXlfR/FGO4ceQIMWV8XpUr2NmXTzic/XgrmFEVXpMu
PzIMcPyzvtrx+goqxqMDHjW8MlHir4ytT4aJlhFyyc+bwCP01TyByJbdCgYefdrd
O185z3DgLpjmXIY85ICA8YxQHgosnKp6ZdHJtZ7RubQoAUj4vRqtLl3KUcIMYr9L
x+9QRurg2LzMeKC+ebdiUauzP22uLDlXiLjLmmkpY65SzSuxjv3RDsGpkjrx5Z8i
bn++rg6T5Lq+ZS4diPgs0MB2ezQm9hlFM9FoOzbJVQOHJItj567EB7PGOB7bQoDg
ftIHYIdplooZxh0m43kYmbG7Sp+Eaq4ceIzzL5cSFahF+E/YeA/WBvznEOs+NB9t
kyEMVhbmzijeNpkpY6SZTx/r05jW+6/LflXQCKAMfHvNPAzMYTMPJZ0j8s6fKPTH
qcDzptodLTmKcSjdKbqPeGcNpAKNI6fNSsXwDeQNwmqZkEOsZXY2CzhNfv3erhgV
0Jy+AUJPCLNEQ4jC958pj2Neu9dN4dzeq1uWK/P2g4UNgd0AfcrBI+R3LxQ8a57O
cWXSZ+uK+j+Uf7d6+a7xHN9E+KIU0TrLcIPV+gT7Fz7ppkFWXdVJ2Bj6gk9/wQEk
c9yJeD3nFo7IOPh3a6oa6HCWsraMHLsoj7havd0HONFb2YBNaqTum+2TtY7XwzEG
x4q1foCw0m2wIw6zjXA8tAlmB7BeQB73BTXDIfb/RklT9lk4CPTxm01vOAT9AjDX
dea6r3mW56u9xMp277evHWJn+32oUjIkZ8PBZQS+ZJkD4qawmPrQsVwgpuKbfssQ
TqVMp9JpwcxyXZUojF9k1lDGqxB7hq+yVw1UviZPjJM0gPaoe9Nz0+/oDZKImuzd
9RMXKczH39FTTiNqm94dHq0IywIfmxLDvdjgCAxV6RuR+kNZOAdyskWgjYQvyNSp
3DTeay2BFIPyW0tNSplkF8Y9DFnGhD8kbUFNGdNYD91gySi1bEH7jrBSs7xOS50z
hvTaChegcB2NBBRF9nXodFLmPMrZZ6EsYBEMPTB5LMK49k7ZEMYIoVcqf7dYIUbB
5sMtZRci+fKhXUzv3chxAgiiQyolZVjPjuWKpKYCnJiHFU/mt/fc87Ubta/FPgnw
AZGFs9etZ+rAl6/MO6z2ez/Jz+zsoUzgWs2t7w7iWdf1cR8J2/5yKToffNrDSw/C
80CQRkbZ7FP6RW0rvu0oIPKia/UNCENTAuegrYJ/mo+NIqHN5Bq3GopR7gSH1EV+
Ph2lxeHu05ulY6VfjuNd0wlxG4B9taTP+yqsHjyC4qhlyHYKRJBLMEfUpc1+I1IA
m7jMHgWzJzcTA1FiTr/smIvIxe6Cv2AXT+gPRVmSjLSmAZ59CL2jI/cym0fm5ZY4
7fOgAK58fsc+9fFpFmzOZ7U2SMTA1fyB2AzHrHTasOd3/4YtTpF/uAzM7coUjs/o
dN0f3HgfXWSnWDna+TZfbQ==
`protect END_PROTECTED
