`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
His8T3M8GMgvDSWQ2q+QynuN24hDOsHeFCATpE+JsF+P0KxZTPlZdTqAlhp+mljv
hDTfR2rTFquVu0EkrNpxLw0nW/OzW3MQSQx/t9aQcws95CQQloOmhnyYqb+cjSiy
tdRrPP0BlQ2Av7kE5zZOPCAgqkf22ulrrfyVwGXuA/6TXlvDMWReZ3ZaJMSqnFGl
Dllgvn7w8znxU07ul/SQw2UO2qXA99QXme3ct+rJEahhQgLhzeFKYGgf0YVck79Y
7MDVpMmi67R3oWJqHbcjTbDLTpM05H0DZx8+12qaNMNebVYDcq6owqH+2qyltOMc
jGQW3FGlVJLHdTOQLod1lKwSiRdIQKwl6etBPcYDEI3c/7h23N2yjFAKFZ34w7px
oRKU/5iYxtcBFF1XyY59H8IHotmGYNDavOZnqQGP2DWb7+6+JhSAB1pKZfNBxyja
RGIUqaf5nvXTbmeSsqkReDkL5dY+IbjILp7Gpq8oGRhJSR+0g+P8tdAFWlZqhyYV
9jkL9HAc1F77aGXFGXWvZu5Xu9INMimHYe0/YqfwcuhKMtbSVONc2DWB6pHfj/nD
f/eZU1zmDRIXgUPvleZbbb8AAfQTBiynBrYCHfaCrMkrW/0NDrjYzAKkDBJW2hwF
Ub1f2rbCrpazGW9omYw80g==
`protect END_PROTECTED
