`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XgW2qI/asNiDw2cA+njGIUQo9Zst3+l9QLXOICU94djJt09hkgMSaFu8LtHNLRKU
JR+b7XXTjPmog/Q1NHTxkSbiHQsV9edHDoDiK/aE87+p9BSRU78smWYJJm/947A1
2JriRlisVZsAp43nLzMIYaoP9PjuIsn8sXEOw94dnMatLWXZJ24xwxqgwTGFnAyK
rHCPUfjhFFH6vlvxGyedO6mHKLXf0QMGmdhlmsyrzuEGfogCa7VVvPdHP4buZAcG
`protect END_PROTECTED
