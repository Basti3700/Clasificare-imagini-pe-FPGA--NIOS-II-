`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47rF7gnyd6X8ijphUBcOF4dYAAlkiCQXBSzD45t9pjrwVuZHWgacWb1gSk4Cq+Ww
HQgkI3Exrnm4Dzr3ZjiA983AxUezDXSoqVt3GZriYAV4trBFAKJkIl8xyFi5omPV
78SsSccfdG2b2SZe+OqOQVgbP79WjXgJeol+9fNpV8Y5I4NrkqX6B3U/QtDFliSU
jx0QAbht05JbFIGr6JxA4No8Op6l7lVpJkQqQGxuBw6+MVkcoUvPYwrziCdcbEfW
3jfLS0QhetsGw0juMTyHUa4O+pwTEwG/TKsrrnbrUefRjoBL86wooN0Y9FTJ/41B
VROJ3ZkVeCK+iVaJfDcP00KKyDOnMN4NJZf0wx2nSu2UNdT3cxY48kncWPXRGAPJ
m5Vn0k80NMW31EPsxHqju70W0lAc1aWNhOwu3Eyhcz8MgLukYxaKJvTy5z3ROjZG
OCY8xX8IhCPorCwVpGbA+g+4++JEcMreXYaO7glvg20Z3XjbQfGLqEg4llWOmfHx
2Wom0QTJ7T0otPO+DfW048yXAqDM0D4v98acBlPnAxeAlvNcnHA3O+Qwa4Z6ie1i
Jbz1JWg3ZU+5GSlIAXNbWA==
`protect END_PROTECTED
