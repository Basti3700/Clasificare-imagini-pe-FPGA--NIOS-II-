`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubS/4K+dA89KTIwJDISeIe3HtOOCeXgXQw7cO2PLaGLqGZIUoYqyqrBjeqmTenU3
CWvOp982cbG6K2aJb8nb+8iPSHi0jKXlV9Z6KJklstNR4EPkEBM4mGvcGadLX8/f
GUh7LAhxdhDE7TaP1X3Na2MqTDIuNwp5TQuHqqZcsaHWSxHrEW2gwTe7jBg3XFQs
B/zNByw6oFTq0VEUc/OTbfORp2pYViUxEeLfpeB7OdJUSSWO5i+NM0MWyFV9Zz46
`protect END_PROTECTED
