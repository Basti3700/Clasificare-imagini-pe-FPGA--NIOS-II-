`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lrrJJvKe7xh7zyKYRNTf2R3MgLIKOwZqpRKysFxDL8/u7FK6/7FPJ+/CHf03W2dZ
OBcZT1ZfySq6r/OczwAdwEZiaOKA60uMCZ3Zm3sXO9A+ae03CrX+UnOVeLRv1Ksh
dhmde9LNdiKYPdsrtUXxvq+c+2KEtgzJ+8T0R4qsDzhmAuWpXXQP4vQG0r2uPWeg
GSrx5SIo+fmXxCly0BJkYgeYw95nuQBrws5KV24jHlA=
`protect END_PROTECTED
