library verilog;
use verilog.vl_types.all;
entity altlvds_rx is
    generic(
        number_of_channels: integer := 1;
        deserialization_factor: integer := 4;
        registered_output: string  := "ON";
        inclock_period  : integer := 10000;
        cds_mode        : string  := "UNUSED";
        intended_device_family: string  := "Stratix";
        input_data_rate : integer := 0;
        inclock_data_alignment: string  := "UNUSED";
        registered_data_align_input: string  := "ON";
        common_rx_tx_pll: string  := "ON";
        enable_dpa_mode : string  := "OFF";
        enable_dpa_calibration: string  := "ON";
        enable_dpa_pll_calibration: string  := "OFF";
        enable_dpa_fifo : string  := "ON";
        use_dpll_rawperror: string  := "OFF";
        use_coreclock_input: string  := "OFF";
        dpll_lock_count : integer := 0;
        dpll_lock_window: integer := 0;
        outclock_resource: string  := "AUTO";
        lose_lock_on_one_change: string  := "OFF";
        reset_fifo_at_first_lock: string  := "ON";
        use_external_pll: string  := "OFF";
        implement_in_les: string  := "OFF";
        buffer_implementation: string  := "RAM";
        port_rx_data_align: string  := "PORT_CONNECTIVITY";
        port_rx_channel_data_align: string  := "PORT_CONNECTIVITY";
        pll_operation_mode: string  := "NORMAL";
        x_on_bitslip    : string  := "ON";
        use_no_phase_shift: string  := "ON";
        rx_align_data_reg: string  := "RISING_EDGE";
        inclock_phase_shift: integer := 0;
        enable_soft_cdr_mode: string  := "OFF";
        sim_dpa_output_clock_phase_shift: integer := 0;
        sim_dpa_is_negative_ppm_drift: string  := "OFF";
        sim_dpa_net_ppm_variation: integer := 0;
        enable_dpa_align_to_rising_edge_only: string  := "OFF";
        enable_dpa_initial_phase_selection: string  := "OFF";
        dpa_initial_phase_value: integer := 0;
        pll_self_reset_on_loss_lock: string  := "OFF";
        refclk_frequency: string  := "UNUSED";
        enable_clock_pin_mode: string  := "UNUSED";
        data_rate       : string  := "UNUSED";
        lpm_hint        : string  := "UNUSED";
        lpm_type        : string  := "altlvds_rx";
        lvds_rx_reg_setting: string  := "ON";
        clk_src_is_pll  : string  := "off"
    );
    port(
        rx_in           : in     vl_logic_vector;
        rx_inclock      : in     vl_logic;
        rx_syncclock    : in     vl_logic;
        rx_dpaclock     : in     vl_logic;
        rx_readclock    : in     vl_logic;
        rx_enable       : in     vl_logic;
        rx_deskew       : in     vl_logic;
        rx_pll_enable   : in     vl_logic;
        rx_data_align   : in     vl_logic;
        rx_data_align_reset: in     vl_logic;
        rx_reset        : in     vl_logic_vector;
        rx_dpll_reset   : in     vl_logic_vector;
        rx_dpll_hold    : in     vl_logic_vector;
        rx_dpll_enable  : in     vl_logic_vector;
        rx_fifo_reset   : in     vl_logic_vector;
        rx_channel_data_align: in     vl_logic_vector;
        rx_cda_reset    : in     vl_logic_vector;
        rx_coreclk      : in     vl_logic_vector;
        pll_areset      : in     vl_logic;
        pll_phasedone   : in     vl_logic;
        dpa_pll_recal   : in     vl_logic;
        rx_dpa_lock_reset: in     vl_logic_vector;
        rx_out          : out    vl_logic_vector;
        rx_outclock     : out    vl_logic;
        rx_locked       : out    vl_logic;
        rx_dpa_locked   : out    vl_logic_vector;
        rx_cda_max      : out    vl_logic_vector;
        rx_divfwdclk    : out    vl_logic_vector;
        pll_phasestep   : out    vl_logic;
        pll_phaseupdown : out    vl_logic;
        pll_phasecounterselect: out    vl_logic_vector(3 downto 0);
        pll_scanclk     : out    vl_logic;
        dpa_pll_cal_busy: out    vl_logic;
        rx_data_reset   : in     vl_logic
    );
end altlvds_rx;
