`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6QLb/i8dWSx9pLJUvycjkVEjJ8dOkev9S1neRjxh+NaasIY9JyEnc7kSQpgg1tf
3CpslEfEzPGUKwWPSSDjzxlLhBXe0E0IOYUwYxhegXcZhjAFclcW/1w35WA6QfQa
MDwCbEo5FOW2fa9cJ3Ai0ifQrAaG241KxdKc9VWpRWEe//+ypkpBWcVe3gRrQy3g
/m8d4VLJ7/iVWqZvczDCpGQtxMiplcpzcSyI7ifLxjMiDD+aPM0/18OjFE52x16+
qctA2l/gDqGUxOeltGZ/Dekel/yjyEonP7ydJDU0SRsBrd6q8y64ii7RuxZ5A9Ab
7/h+9l+Ei75eEFS8ZkbDzHi0by+tBOiTx9FXG4XzPbONUbpJwTu0AGZoBtBqWWei
VqCttuwMQbvr7XmPlDUTp4oXzjPRtX3t8RhjIxGCfRufmXNcmZSrOm4c8zIsAunl
S739D2dwrouCwtRdVwXqcTwY8M1oh9i5Ac0p31/fCrl+cHqeO0JQhNU2147fctNr
rzorFAMiBkUmLva91ktoRJtIyjHF/AmZQCKrpRCAwkpm5Nl4N/u8G0dAdBKlXKYE
aNNQw+fTpQ4SmzS+NkAWYdtLqjZC2k9dwrqXSrBTg9Wgy74j+1l/PoByOFnLIOWl
MnXY1Df0Fhh4I69WLtm4VCBG+Q0jCk0xt0WusIvtG70=
`protect END_PROTECTED
