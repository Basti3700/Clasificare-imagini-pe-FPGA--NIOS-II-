`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ikYfhxmn9SQUkQkY7SpyIrEE4EJRcvPe8pKB7H7e+sd5TG9MHR9ptKnBrT0tGGJo
4wsRlFhSV4xAid78IlThjjT69dqaUe6FqVPuOpzX/IzaAUwLIyciSU9SCQNluZkd
m4GRpAaK//ZD7W4j3jCGd7gdrqOWR96VUdlDeadM+zIye/vCX+tPvh+9YzslfGBf
Rd+zCg0iNJBBPkLuIXMGryuvDplDEHS8P/RANLTbvzM8lY4o7DB+3EqmqfgGrUu6
REOL8Etfj9CHfbiskE/WMUKdHrlqfrZ600+axJ6MoPMMhkMan2TcTRhP9pX67osT
A4kLEgjpJqW1n1EfOOVoVDWfERQHr9lFj/K6j8E1W9mhrXpIDinW0sEPzK++IBbG
wBdj6Clod1Qfe5C0pLXm63fgd12XFux3J9g1TeiMa4i4kRxAO11cMIqg0WwdyAmm
d/zkZDlx/Tt7kgJ7LATUMOIiOGNjptybn0Wk34nOBtYR37CdPUpT2O3cDm3pfTJa
WlQbBsacKboXVxSSX8G+KyHDiMGoEz9clxDoOQQCfbtFLiTvzDmB816NeDLdYj8m
eoZLeb3vhaSL7Cl3LJprN0jAl5N6M3arEfbaEYdOzHuojz2J4jwV8KT02LA91iIU
B87POU8kiMnt61t11lozmGLqq9h1R6BHpL3rRRT0LaI=
`protect END_PROTECTED
