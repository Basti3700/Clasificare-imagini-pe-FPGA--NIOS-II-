`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDhhssS+8d0Hw0JGGRH94vJzC7kGMKnwQkV3fdSN+iC0rVUMgoW0KQaPmg40cVwu
GCsy90Y7e5nxGiWyvQgipzYp7pRMf2b3JKF8GB6WRgXvHp9p2r7Jh4ch86aIs1lY
NlV8NfPciI/uZTHhKFMPOZT7cAIdgjKBA/rXyedLkHQ5ON8g2WXDFfXivNLzUMyb
fwNF3lXJ0lRxsHy/sqx4U/O1kmRt5kODgcc65IBwnghV/XiOsT/sGOuC1nBHlgQ5
ZadOccxfu83XcD9RAqslKTJlUF21+qnPszkQF5uTuHsQVlccSy5JmysgNvzg7qJn
aHuzrdXuC21CNU4iPGbxs50leCQ0iHTUjF/bsvXDlgnESZPS9qLFFBDfkNUCerE8
RvckJytWo3lDXd/9c7dKwI9w3Sr5Xlk3AGf0TQDcfUrgISIO80+iCg3PrzI+FrE6
8oYyEjMWYMwIbL0fHNj32FE/blRsUdK7f3F5ShsrFXrJgHP/0h5Dr7biXo6jD8+Y
AokCuTiajcOCRINafWgOHg4TAJDZK4pb/SbicZeZ0Urstwzx2Ji/MBDGCa3huxhA
dQBNTWR0cc/uP5HRDvUZz1OCFNPonBkkPDZN/eC0O9EDWpEoewqe3DAuxmaJycxx
J0dZg1hC+MU1DxgCnTxyLLrCjvAOeueGNMWW3MHvupLECUXYWuTrfzIwKG9V5uoV
4NtR6HsywsZLFXQa57/W0w==
`protect END_PROTECTED
