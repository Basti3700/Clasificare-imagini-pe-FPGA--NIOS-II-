`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WOnpZkRZ6Im0pKwe8RG1QF6e8oOeftfO4ueB8w72EIPWVv1MZzp+7arjWET9Tphs
HtPhFEDFx+Ss4fiGGdVO4RHFyen7p09AXvZ0bEVm6iM5+7jGQaZbFzfkPsVk+WoN
4FGhlU8a8mrl5/X9BjRRjeh+ZywI9uh+MSL2x06EzL1cBxhZjZh6eS9qbNDHKY7e
Gaw1QsnvrxZ34oWB8OhW1o5Ea5KZuljh1PMpirUhdrH1ZnHssvlKJec1SzIm6Q4/
fzyn2Qj5paWT063xzef6+uLn7kagMaeQnf5D6uhRB8flrBNt0IzEZQNWEHlZnu8j
BF99pnoE7H39GGNFXAhee35V4hBby1wNb7wrcY2TlvvSKF9xjylxnmbzsltowj9O
BLSnko3r+gi84P6BRhGr6sNkjhQpu3RbMJj3JGsAIlj4LMueMwXBir28jW1x6aFr
mVcKqDT4stNOG5V9sMY+IAfZp6raTpDSSBqOJBpJXVXOaa3B4DjbdjLOCjHY7y40
Mn0lGNs8rDSfL2uhjfacS81Hk2dsv5WF3Rd5yCvOFQQIHbUmkVaoIyK1nUiAzt6g
QXFfNSe+pZ/fPA2NlYb6HDRAC2+j3sHURg0+d4QS0AZpc2NUsngy3qpkOAyCKmQv
rBIIM/f3RfkmsewOJc++gTL19vQ3P9vH1CZbL+I1IMRfOl5KHZ+92EkUtoCqPY2o
s5JKoNlYA3YTTdjEK/d6dUbcqQUReB3tYOVYErVj89qScH7ud82rgFcXmiNrfHpN
vaLy63QGXC0cCmPqJwr5xnCAsu/hEacimpqbUsdR7Bc=
`protect END_PROTECTED
