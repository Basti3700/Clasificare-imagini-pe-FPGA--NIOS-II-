`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cdzCi1gZEhBFp1HUOhzhjHbb0cpBNfasHup++m9vupiRkj/v3CeRUwhEbCqw0Sz
AG5ORSaWM5nCX51fEHbeXNZm5Oy9TmzdH8jAEjT+mxg583rk8V+RJ1pGwYq63sPI
je6w1uWYha7bovFpLM+0vuS9/diAaOpZvlgMufhKmbT619zII2rDabEemD0rlsHh
9ZJUlO7+5O/h/58q35WkUrnBw6YEVpk9cO+mQCmgw+p5/64xaigAtcL92dB5Glmv
qSqMfTjXIfXFa2odS0/a7f8x12KNkWCL8Yl276+JOUb/so7JTqrpTNiliQs9amZD
Zl0ddBrtiYoJ5+wQGw8DJ2NndSgCXaY+NRctQP/ni3blk0//zzVGA+aCOsehhHuP
3y998WKiZYJkl9r3ONMPuhcDSXgjiUkHVnem2c0FcDP68IWcvwr4ih7ho7PDnJ4Z
bEorWdbRuddYJQSy/ce725Q1rD8LunZqLBFJUDpttZvYlC/75FHwr1jxKsdYOGg/
r7xKPJzYm03FyFSHCYV4av/Hy3PTa3M7VpTNc78SM4ygfSJl6YtlTolKwPqPnuE7
dDDATs+f4U6hP7EtZREqlnRe2zE2Hat7bJrZJpq++YUSRr/9CaIgEtfNY54Ci8Jm
jBi1IZ9qQliRWHeEEcDAMJSBagzPOJkuHjXr1q1s/LKtduRJPD3FGip+M8YVyjBh
k4hNFr21CYMFwSHf+JdJzx7FV8/3tRvLsCaMlY+8//XDbv1acIwycDaw4uCqx4VW
KNovbZg+3f44rA7iierQwp0ucq2gJD0AGysi8AYCbuajCHgXFIN8TyJ47xvwZq88
zbdRimIzuUgXNGR1RaRL0En04XvldClSFRz+qyS82mEUDsWBp1iAokqiDM/jfGPR
HbyL1IAXBIOIyvbvuhoBTeHROQs2Sgrk+n1YnS3EVoCARecY06g0qQEOXGJd6D0L
q6jAIVWleYZ+RJwDfj92CtzjLMap/AAHIsgRIEWzn9iqbwi/fFOdKl+VwMiGVoSb
N+Ac2CyHfpCW0byYs5tL42tv9DOwzYAXBkOZvJMxAr4FZqKsV7NFDjCR6PITStog
vRrexsOCmCIZI6sAiBKm7z0lATbwYnbpzrX468s+4kLbWnLWHVbq/NEOzGV1Qgrx
6L4TabFs3+lW6ZD5IgCTvrIgq5EuuXtNmkQoY7Gdpov/HdCT/4JMYg6AZI2IMo7N
+rx3kDrgRCw7CaldkdZey80r3cbA/Aic35IlMRWU98T0Y1WwT4e+30V0t/KYlcDR
cXEC314sbQ1+eWyI1xUKCtyiStgdoD6VvL5zz5pG93aQu+y+ZwrG7MeZhL1NA/Sf
+AcZxLQ5TcuDjdTo0ONQTFjmcCEUtxzxFszoGuIFtlqQdNw+IXK+ivKALaY8iiEN
encl33u11NbroCoIGFZIuGoZlUP32EkjrXqu+GkwZu7Hj61ymvvxARg9Oh+FnHxH
S+OjhiA6JJA2AHMQGUX1srcAAfm2hw40PA4cQIgDawK58tiO95H+L//AsXMgHZAS
F49rPn5e8mM+wP2Ejoe+6Cy3wsV2nOiYT+DY6+sO9QD30cadfDu2dgGLWbxqykKw
D1y1oTKXWkZ0Gw8GbuWp7U6n/jgNCMhSIanRHO+CuFjB5FJiv+hdSO6WH8S0sdYn
owq/A+U55+cZMOzbpCMESLPcI5sEbVoqipy1qWZNkC94zuIJtVY+BsDJcRWAo3m5
O9G5gisXyJ871jCSNyEBq4PjnFEtVjhvDWARy+cHjzP7kMFUNMpq95RYiMziSSj+
+FZnbz4fnSnPuRFQy9mHibeebAf3lYGSpkhkq6d5lddYsiZ1looP5Gp8mxomota4
HwtXGKaAlwDy+97+b3JqP1M6cQjj0mjvnfKJ6KhdlPs4bZxWGIAEzNlRTzUdQI3q
7umVSJhYO7MJN7jh+Y/66BIW0ds2gpkbr/iF09ExPWRR+U+sFqEORCtWzMvCzxBS
CZ0i1zQoas55YKTmSi+hA0fMWQYcx4hXlnlXbA6lj7pDarvXXrpl8+PgQrghr0Tr
LFRUcvEVnI6NGgtie2wiu/QETbhlxPvq6f2UH1cWRJ+yxIOIza65lTE4e50/4o14
mcfs91dZctnUWxDe9Bmo1MX0tBlIkiKSzwhqT7SaPrUkzLu3H3SbLytT4oipEiLl
5x6l6aXoyFAnHUAcGj3aWESUtH22/rfiFFlImevQnBcs+ai2wXOsCSgHH4oLeASF
lwMdEiciFHzb15zET3kIcmsqGRSe28tSddyJfe76bYE4tzzSHc/u5ubcgaM39nSn
ccbXXROAtPXc9fzZnMGTRvhksuO1Q5EuzBSy/4FYqSCFWSJS9ydXf4XTEY8S73Jq
MEmeDfNLWy20oqeUvXBddvQ6EnFZoQGpi150qpZ+7udY/YS6125AalSKaR4QOuh+
TcFn4N1/hrR6nysRjFcwuEIWfzF4PfxvGphEl63raNTVw5Wu/7/bnApDnMhizy+r
kvNiqr1ZnjYG7nZ9MLtIbCAHTVbip0o5rJ4qgJH+gkr0VzWTjCbXEk+/qLYUK5Hk
M4bcHpUWzHwEfMTx5hYbcMd2RXCc8LYlpGRR/FxPvY5FLFy3F+0u70eBgzO8phk5
fVd8E7PYjhuz7Y9YFj06LsqlTJtmMwUZcaYz4Dam3UIKtNxyGcgEn9uoXG1nAwjq
7xP5oyPY093BcHZ+1m0Gp52CNgUEIT6HcOhycYA4tG60NrnACJkKwIfA1jm6QuC2
iVdskBjSiioreyc4LW0kGtnWk4aFScozWxbVJTlint7PboKHd7sOOtGqB1AyYku5
AYx3bKsiPmxCYzSuIAzklykdN/0odBLfRUufJL9rS9hHc+KnpjbLXwXkWAcwei4G
/RmcIuFfEmRW9o5j8N0p4Hzu6K0pqX6i3Cjyg2YvKosoLlqviaY/p7aqRerdC3Yw
56/NEfjZeXnPn/zeofxt3jJSdwrQmgRZtX1edvmcgbTMMH0/NCBePRLOt5qV16Ff
oUMXm0o4VukgCU8ib0xtdiqwwEIT4IHRF+DTU0HCpEhV+oaD5dgvROdxOVbtmuNS
RDNTfn7g8FQhBvn4Q0aSzsnPG0RXnlVHsBUUyAWcCB8mOz0MsLvOrn/3p9z/b/8u
xJbt3xox850i+C6wPSF7SbcwLkRYwiSFSUTy1yutAYHNbCHcNzakRqUgtpyLTdDg
E5jzFowRTKtgLTIq9pzmrH7pejT2GBGc9I+zyMr3mXoPb1Iao0TkEBQpN3S8GFTJ
iz0QG8QG2LuAV72f6OZ6ISIrpUORDNpR4v0h2v1I1WiqQlv3PeoJPTWPoPlVvUIh
OEdfFlTZRkXA6gDTL1YhOhcrJdMXA16H8myFI/KvazPaVRiDE9icv/0nflee7F7+
iVxPk1q2T5EWLujm96F4yAY5/Llqfh5xFezSfxRv3d+eFNMIM9Sn1GfHTCU76rzj
fvBCKagBD3GtZbGx3g4fvaGb5L7V6moilAVuMIzh8zHHQMujBcrIJBvEoxpF4lJF
s1Xvg/quxGoQfazbPRgYzVRJLpx3UhnSEVyLbU0A2bEewd58imnmnrSffvqInY06
TOP/+nkjwhXshq+FH3RpzxgWwtBaoWDEHO6TuQ7Efgdgfx5v7CkDesHgiqpdUiAM
HinCZTM7ydu5tDbJcueZWXlF4lU6CZOgIn0uvJY5m7rJpUhq5TZLBcgiU3XLp90P
ZkAgOK0M5RU5sCLhwhBp5XZr9oQ0DML0U3OnCIv1MynGtNEY07URKuOjjXr8ZlbE
Z9L/VZNVr6PtsJm5MNv3oJ7PQeVduXcn0eXvB5LIBOfhF+c4wZNTky+Z4gcBuVOW
WY/2Ta2MKdmtRn/liiGG7FZKpbrRpHDUZ0qe7gVBk2zIyYjODIG8g8vLBmQ0wPlf
SDUWBRMHTw4FNm0W8Ufw0Q==
`protect END_PROTECTED
