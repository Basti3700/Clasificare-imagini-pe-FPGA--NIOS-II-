`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZpY5aqoCZGy2qLD4orfU8Z3IRYvWtdXD9pNXuIJlmf1OzWZ8IuYSr/hS1yYD/pX
LIMGhnCBYJgWQ7XgaqHJvf5aBhUP/Ko6Gham7YkZ2PnxZHd3fdlhchlCwSL1Jz7Y
fxc9EFoqI8wAZ6mjiRIWkwahEsu/4pOllG9gwfdBPT0zK/0AZqf1GqxKYmqK/OGm
V3FagqpkuRelHmABnwe647am9rByT7WE2jHi6XXQQMLLzXnar0Ei/B1whHsynVNy
YKPkRKCXr6ko6DIhZ9l0+j1BSoFGeYyvoH6NXh842IyXGH4XDm2JlOkf/v48l5tQ
HMMM5utNoxqNQc2kuNGwdAYt//7OAEKXHDQ02R6nzPFp76OpFJmKPf3Ze3DJIgyr
oomgG+BHc/RW+rz8M8DD2H9B1ql26ighey1acmJt9KbGtL+k5tSIU/e+X0YvZ1RD
pHpJauPRl7E5Vww/ZGkIIC6sfAl8KYsKd01yEYxaLO1FiyGcCwWsemdEA6wiFtz5
`protect END_PROTECTED
