`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fThRG8MHYY2FkpkypUryuLAZ/zoLqsFOJ69nZ2KPDZm0So95Mvp1SCaj3HJYc3nD
7ONXNofMjMVVdj+K5YP3tX2D3olOmv1iOKKM0F3RMifzHq1FcopaD3DsKB+4hZ/Q
AnxvcgIUSFbUxYwrF7ihtBpn+UmNbuzCDAnXR5bZt8QkBqXcwYRVLNP2zIKxXL9x
9uWk916SFlwMfzCaUqz+hXRzutZ03nf26yW8EKqclYDLhnRKMK9HCRFEAY+8v4pX
PTUzoWjluTxCaY0HKUprm2ReAFUWGPiD7I/eUHWRYCwDaVLp2ZY12bSQDyFVFe6D
8q8nLMLvZyEIGjqLnH7Iao3TDcX++LxoT4l8TWND4wfV6dsxM4UYPqa/mcVmvdUq
D2o0LdWKaM82oe8FkAgUAldMUdiVUohOzZBo2g7aBGvxCZReSjtu2sOSG9FSu3v/
F3aYKHlP0902sksej0oIpMuRYoC3PsxHiDk0VgVQooRlRedx70tG9U5Fa3Xb5I/j
a4tg9Vy8oY9ryXQz/GoXxiPmuBOnZer2zxzDFCoEfasl9haISw+tyz3ud7PHWZsC
twDIXpdIgZ1f1//DVnmQHUxSuyRcUM/0WTsY8kNoTOd7wUoZ+xTX5XT1GYQrkcvv
lQSQqvsmeDanMuRBov29Eld1vwRA3QL85hW58jYvkWMuuPNcVFUE1+mS1dCpnHoe
PVRZ+WvO5bzotk0TYA8nsM6Uu5uUA7T4Yf/nt/4EexVfwyme8nOe0stmhRbdVfXq
TqeiEkzb3hQwB1MiEAa9bNMog4Xw/HqtMXHtBpOtMsEkN4uFHYsWa9d742VK2DNG
s5xYUoVfvQSZS7sfbSVS7GqzXph8qTq3r11hiPN5U1m5sWamdIUBYWHflSZGdQG2
4qg6AkkUQBi6IVU7E9oLI5R0i8ShWmgDa7XotXB+Tyha+VK21wVAxBTxeHfQuFD1
Jg8VvCgtD/icH06M057wgYsV2q1kUoXIBY1PjXjrFglwoxH+vlECYJRmT2reYles
AZPe/mVUFCIGl3A7OQlNPa0jgncq+kwV4D58HiEAArv6kiGNKhdp3RH0Qh4FCt0i
1sPhiXZloOPvJWHN8q/HyRGCLWT7gnjjk7XKD+rCl1HwO1kB3f7xQyViF4BmyM+h
E5n2qVzwVRw+CTHCX6Ecd5S9kjk7uyOdb9u5wV5rieq9va+87EZmvyWCZdHhSkwB
DXf75h8WXw9BElQ2tfJauNczuROoX9d5BKHCsQNq1Uz6SD+a0fgu/58QydSzRhb8
78u07Ja7LYkoTslQSffzDuk7EH8qMev+TzJ1WmiTd43f+ybx7zDMVyjiTNB/HRkS
LYzdj1KuqUOVsxyYfEfqvHGze/3S8kkAsJC7xHULE/6nBXhbYYWUOGZx53Ir8wlB
mYfuwsCN0NWZpOPY72ZNPnJ7hK8qL//GbeoBCCcT1PTULfiMPenQaDtpTHnUrVqf
vXmP+IQW1M9zb5TN+cDJmZdxPh7RLxkzc8k1oySR6JPknruziF6wdCeqPTXaFhdP
LK6DDReDXom2N1ZvZpk8Opydnj94O2l/Qp9xCHu4Yc0TR6kq5msMY28DFRkkVWvP
SIfpZKIeKNcl6MZ8F4+pLRB2GVkg3lHwONmx1rFUiQ8XP6rgTHArA3olLQQ0m0wU
oW/BJZ8LIur2etgd1WQ8UkMQToibP4/8q958YDYdVk4iSE4IbE5PKS4KMIwYlNyK
HLikDmywQ6QlzqggGIrG5g9oBtT86Z/ZYGmxWW6a4z2tfvhkq7hJUSMGMPAjv1Le
OWPup5pG07mTtjpBbgs6FtA7GaPXnySsR5KZVcTeRkKiS4Si8QOs49RpXebaaQsL
XfckHwcLWNisjsahtXvfy9bT4QFHZpEL0Cgec4rGmgdBQZ+ASVBwNRT+Mh3CQ896
dGmc8G6ISV58iI/sQj07C29b/FbnVBOj+p8Zw871aiTpASW4PKhx8XKloaYDNhvO
GfG5FBSxBgbp+SaAvvjjX76lObL19RpvEMGsd9mBbGLCGXBlk9sEO1tffOB5XqYf
jeJ15dL/8wpWxOw4+/eAk7gLTOdbtfLj2ekDH/NPGcg5TZ5hoO2PY9+9VloOkyfV
CV+ZaR4U2Q1jfKapiO24De48hMqDQJqfm2a7filcn/R/0DEcAINo04i3fMOm9cl8
p+TzPApppK5eysXQOpoay/oE3K/xpgp9yCd4QAx6hRmOlbhvc7fAAv6pN1kChS5j
IaNtJCmoVze1at0xmbLVHKUVnOB0sZmdKhbfyDN3u7MhGjVmO88cCFspBmb3z2p8
x7NqjHTh9e155HmclBRZTUl4yeFL7l/tjoTUd9neG6UQQbIPiBn0X8375u2YbRPr
`protect END_PROTECTED
