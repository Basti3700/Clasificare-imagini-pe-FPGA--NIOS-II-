`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
07u1iiH5pt1ewZJ4c1s42J2vkAzVthgylr3o5XMaG6iKQsy3akYdklufukZBKJ1n
ygbxm2F/hBtm485+0tiNt0IQnwdzFPNcb3F6srbu82euVshFxGI768GJ+9RMWjC6
7aulw3tXnNk2RGQPqG9bEz7zUYLFREMveyPgZ3vzVCtzDvHums4+MGfDoGdbFWJZ
wJYUihRWRDos4XfXosDuvKvy8DLAD7kYLRLJLMMTt1d7Fj/hhFEwEakKUTJP8T4H
q7J5PToZPY6B38bzOLk6m6PV5pQs3gdRT0jaiCS3990SKZD6sebkWhKBcxp2gMyH
Q5t74sBF0yCNPbq/qrmByhtKLVz1nDJ167KwIxZkZ6moPIaS6aDRVfTMJguTrd2Y
gi44VNjYuiWIs9mh6ggWYCBpzcb+I3OeR/6KWNGEFD3KrEXHZtWzB2vEU2AgD1hy
aE7TfnW0dKXaTJwspkvCKxzEt4HtFU8S6Fln+Xe5DZExeFMscRMxNcNrlKk3Rmb8
/JdTQ1WToBRGCgJYKGJDzI0TVwQLjyTzK5Dh5+kSiMprjvN0M9sN2oVogYVZuRZT
J7tVAmgJMDOfHPUS/gwiW41m5pIHQDcWNZxkmRevVsxJDBgv112nhXjV04z1CqLo
6nW/zxGYPNsXpDkiIvqc5i57S00OKhcurwPoTzKuZZrzHXk/zSOd7cWQxAs9Fc7O
1y1mxOGRbZCZHI6eotQqYBBpXa+F+sWVvQDeSQGz6linZRMG8YIU/SeG6bKzfeHr
m4r/lzWc20To2mKsbAtuEeUeVpBgux8mJzidUkqF85mDxsWKXo6r0Zy/95ByNpsX
9ivJoE5a5vp55YYoFxHu3X9OZXBKb+o6vzaGzMAOIq0Pi3tA+zuaKR51W+h/pbq+
vlMjz3mwls7/sF8UOtWv8g5oM7j34ZaM375IiFZMMtMaXvWtfOI1Dn8fdoW/HGSb
v67JFznk8ZRNxoBGHdi0mu6xBP1Hx2T4tfXdeeFKX5gKp0vjgia2E52Uzc9K1Igb
V/54cn3akoKb8l8KBxQ6P9sbJ7kHS2iVPclaAEBY/l/zHpHgYq84rEx0jDa9pAAp
i96zgE5Kzw/lh5I/QAXOl7BvOXPyypXC82HWKFFNEzZRg6WtQ9OUGRNEs+mFLlhG
t1V2u8m4oXjF6Y4y2M6Qz7MW1sWzM5i4tWYrOD2/wssW4ZhA365XEj2lZhRuotOJ
xtYgB99i9CTc7WN0MY3a3Befsg2DyI5k+cYjUkBw5mlz8ZQtKsYCiP2IJZilRa6L
qv96l4POIbXTkN4bA/TPW7eqe393TZW8Eb5J2JPdQLreFRMB5pXrCRrcl7WYqV6o
NGhDH16eCAuO4YguIDvkNCrDiImuQpbU+/cEPNuZNcQ20d14utVpf1HBEUrN//V3
yWm5m8JlS7oVvbkY+yd+HtUqnT0Rgt9RuyUieYxeplwr7awzzCJ8ajR2pL7gj8Lj
7ZHmNQjFZ9Qq1ugz5rjxxANw4Sq0lz8AD7O8v8EOHI758Ww70vRocw62mOte6tvU
W6++SsxcNE9cX4OY0qAm2/INS7+a59N7PiMRrlWwjPg=
`protect END_PROTECTED
