`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5r1/kPd9fVIjqwSM6T3gRHQkPcNtl124gGOdtDDA0+PEtxAvTU5ugirsd9KmKBgx
mRZabf39aqPJM5QoNU+8CsIeMkofRKiHYjIMcBi3ZmL9UCIm7QI86ZPOAG358Lqa
PBrOdPxWV7F5hVN1BMHikd5Szb6V/lck7nbDW6suoeBS7cFz5iQIFLU+Dbs18GOg
cUUQE9rqsYeibHt9qG0tm7g2XJXiJP+PrhMiIla9OR1iTR/QHHlZxKKDTYM8AWw3
aC5Mkh2A0G5PhGsQlpXprliyYEDvwAbCj+afMpojAgvn5pNCxrmZ1k6wv4HLR8C+
q/gPxta3vecD2RKXNZ2DViUeE6TST/lnFAfBhHyI7Ex7ekJunYniKiJEUzsU+lmQ
`protect END_PROTECTED
