library verilog;
use verilog.vl_types.all;
entity fiftyfivenm_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end fiftyfivenm_routing_wire;
