`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDZ+hnp+oa/lVAq+LqAqN6NfESl94AIVZbDQruuitHIG1XamcJ3kqzg7BSxAwiat
O3qLWzj/SAbSotYFOkXAHUeHxS9BV85sfUyUei3O5geWZX7uQnoKhgRuxIh1FBqE
IGoHq2mnDAFw6Jt0k0LLCqdTNusADDgVvDHndklzMWQf6P0NbBOldrZdxX2as0Ab
qCHFfVdt9b1W5saiijvw2yF54Qf8kIk0UzCr/EwB+O+VByssE5f267dqpaLscOGo
9MiXIMmpv7KAWL6F8ogCcCKDqyhq+SgagcV7TSBvUXI20PbOtMEgytxR4QQXF4yt
OVTQJ3CZJNXqwMPO2hN5aNWfGn0cqEqOcJIET0FTzng6jpJy48o93cV4sWvOFVSp
d1+dfR+udC6XK/AvANMTanVYSbaRdEqeG8hH1MiCXHsj3xvcwOMezqMMFMxKG/MC
6YWhv9+9zcrvbJ02H+lcP8avJVSYnUHZ2SFL7gNg/hGgpVs+m15L2KcrLkTsIIv6
c1xy39ctoD+d94umXzuawshef6zE3EK9V94WT2X0+UGpLX+mypPaCtvszVfpJyEg
P0Fsb104HW+uXy0ht2kgEKVpgcb9fSBM9W35lGwoBAfGJYfHzs2fQ7a26tZYo3jN
xZMbslQrLKotaFsipNzbbE5KpY0J2m73bdsriynnMS4=
`protect END_PROTECTED
