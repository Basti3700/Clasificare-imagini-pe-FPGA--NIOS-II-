`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ub3HgGyKijYncEH1y4OqDqi30g85Xr0VC14aY2gvaXF383AyYRBNbHkSf2SsGBPX
0H+IZOqDxBGKNfh/vlv3pDiUObCHGvxdGLX+121KkArKHLu+kz7+UvQS3RbIjcbs
SiFBLVbKpjDhZTk4WMLGLnzy49qzygb646JfvQ7A4DjQvNv2SAEqIA1IGNKXDRSz
UZ79BrgqEYjzjk//dosbG2ErLUrHfOPWUIozVcpDvEQojMPaUvVGtt8yi/gNYlIA
`protect END_PROTECTED
