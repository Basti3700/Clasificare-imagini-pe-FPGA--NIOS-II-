`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljyvPe38CrL4EO2KsgjuYrrzFY6xxdzEVEr7mBSKBVMj93ApBv0ZdgzhW/eSQylD
HTloDG538UOjFSYVw8UxVfmkM38bN4adQIIZej3EdzdRlixiC0TTbc8DQXJ+N5m1
kfRQpIT0lE193aAlknsnVv5wJ1x4W+y/QQT01wbf3bF03uu8L4nx2I3KiIpYHoSK
zKlbhrmR6Wmptg8mWTow94LWElglDPFZ2ls97cW3HkjT2WYMZeWhWwPyjFgUVHaD
q7hdaVNiyCAGkvngORctwDvpTzKdimtf11Uz87vGbzgGw6LJc++S2Vob0n80zINE
AqrObh0nzzilM8Nm52helzuO+O4m0/LKpch+OcQENo9dwURkz73EZdubvrYMut3O
jw/paejwG2hUCcU+x2TYFTHWael/9HvCIMDNSw27fxW0pnMeAgEnOBTYc7IVcvI9
eAZ75DIDYZHFwlIugeD5SBKX4Jy/LDne4j7oCMetVB6aw5qi05pxgv/c/yRCum0c
CHMH23dlzG4b5IOTQwCc0cpH1yn5Ub9cbFvKgO2X+v16h4drFPHLfDXTKX7+gPBc
w0jfur/t+H9LB4sx1pbKqBhubu/qZH0kF8pBihfg93rPbUFY4AxJufNn8pjRHUH5
aIrS+q/wSEjrfG4mqqgKhCmStpNiUglgj7t+KVQ5N0KpXdkjmYAxpYkWGrzxQtiN
ngo6jpLSXti8YfUcxbltBr4G62gA4HC0KZPZ9nvS89g=
`protect END_PROTECTED
