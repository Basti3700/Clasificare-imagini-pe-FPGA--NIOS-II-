`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f20gdxT2rqAoNRMZKue0mcK5IHZyTqCl70zYdcFGRPOsmFZeGy8g3URgR4+X7/VK
x7vKVo52G0/fwo+fblYycdORku72TBtS9GgQgDu1EAFxIBigjXqXK2wrvxvaP/en
iXrrRaD29xz1D1kKisWAnLJl/g8cNiTP8YQf+oc1mNvAhT20KPcXobPikzwtKthj
HH2ShjUfDLrXmE1oMrhE6SXB2BlWX3udVO7+vQI+Vo4ac7ZhBQdhk9hCnN2GTTbj
PFawgmWeWViWkTMXHXJiCnj07Nr9A/PPNAw5JJBrvpP0yveRR8z21v0eRMYPnLEy
tsQb6WcIAVh/oK3Gh9ZoidInpwa3sTbIk2809KBs0p1aDLwGbx4FJ3L5Pey+JB/Y
roI23ra596fYqMcf1/TeQG4+klhrX6hUsuUD0SiSAOxfuSsWdBmSJPsUJ0jlaTzn
dRRoJz9wWo3Dqic1x1JOAW9j20jXyUEo7k+AUmvaCUE+OnqlTcVYT5GaKnOErBZb
tw8RWGzJ4uGaaNgDPYkxFwXKqO0Rqyu4S7sbuOogbA08/OI0U18pPrCbiAm8cm0h
uUjDiRMGgMDOYfPrwy6UMA==
`protect END_PROTECTED
