`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXmfkui2IV/09M0rFzE9sY0cBT+kIHoqgvWmiXQrIi893O/SghDLZ8nCm6CQOJVG
u5TCrd1Fce3Fm5XaAhOPHBNuL886UVikim+UTQmetplbd0FrvU1RRj8Mxxt3W3dl
6UqwGNYCzbTrbqYJMUEMuOqdX0TcqibMJ+dO06VPBnCfrhLlHkpGUQ9SrrSjvYnP
pi/5RoLCbpSEMwcPjC5J3w679FYcKghVA7n2eaCZniOnkVXKcn6EpNdzeyTegDSF
vob6cgwJHSFlwLpBHXbaNz1pifIJAKr6Ogsikr2KK2WQQu1OdCsdz1JwwHOtZ50m
iIL/i+MEmUtxqujrfMYe9dyDai7WOHHKEvGKqrwUw77RLAc6UosuxIRI7pOvHiRO
8a3+fdmbjw2su/Btl43xQ6GMBtY3rVlwj760RQae7m3HmIqBzsai4m4+Gl6bpAY4
UoU9QPmoICi832QzVXgWdiSqP4jQF/wBrXnl6ZQBR4aKdX4QRsVxu78fkHWgOhwh
SBvVt+u33uiMMvSKd0MmumHCUG8qJBFbxDrN01Q8/EuxU2ZBZcl87TJ3wBhxA2zL
1VLtAFDRvBi8WQctVE0CWcLDSH/U27DjKZFAn+8nF4VJdBaWsHX7x6WU8QCfP6oc
u46LOAvpKxmFapEXnt5fg8AYl5d969wKsJNxFKQwwVzLObJ7j9100WiVokuYwqYZ
oFhAYcPSrOY6A30ZM0ExYU/tQBsziRQTT0+d+6xdSF4ikzr6FjP5ETsZXBd1mhIc
UGgbLuYo0hFLw8KlrHPazUpWH4Bn9qZw7JgeSeVE0hghKNrnd9HYC2+1XdK8EDql
oICHtDgnxmEgI5ZLy5udazy2+AJJrRM06oMOWj+tgTRe8W7AnKJxykPG9l+XB1w3
AXsdaRCbDqypR4t8JPZPiw8DHgPA4v0Klzo1OPHLK0b/2Gb7lZZqlHN+8wYpOWQz
+2w633uWy6nZIRdE5xKSFJMc7YcZZTD4blfS9LCV/7wCZbFiurrH5dZ8h2XDVq+2
Dj5sbHErGoyCnrhjXXo4Xfk5ayEr596wS3gdqGo7hRTvnGnNE5OQYERmlNSPJqt7
BTLeo683f5PqZhViQTO3cybJ/LKnXGryRUY5V6851hC/85diOkNiLxoCa7LUMl0n
Q4KDVVZyvonh2+37Xw4BrRzjRx9E4JpxD8y2z+dJj36EI+DqCCGyBb57na2i8Jfv
tmtkGj5dhAb60Q9BEg9YKRMycN5PqR/q3YqaV8v4cf+h7Uf7dmrSN3Ubv7XUcgpw
6klELwx5DH4w+MY8RTCsUuSV3VCUJaPnGCNr1lPAjVsNUgV6vlrHfAuD5vTvQP/o
LOm7lkuy1frif4D4y5zk3dq4UO+C7hOyj0FWP9UQyIftrZW9P1Ar7i1fjH4ydgCb
qs5CrRLJDQpVNEyVgZvaNhA9j14YMMlpEd4MsI+ONgFrYYPdj0fqxywPhQ+eo+GI
mbPacmVx9XRatK/dPV+ez/G4/RcP+SAKSHhYS8a4gE2SYzvwByebPKcWiTSNuH3n
rDZReKn0ejWCuw1WK4HkQL7rrum3cOxsQ4+lckZOyTBL0mqiyxHJtWYPQlVwtOrP
GrNBXFVb/RCqpfleLGXRXG2nuDew8uP2BE2ZgP8f5GZHzYG2nRlbvJ0G53cBRfMn
rGs6vj2yJVOgeAiAibuzNmp4vbwv+zMWf11DjfWK9lhWcV0ye/n1T/YWvSyf0eMR
X+Bq9WVzMdpIdTHTVTSZm/0Z3Ra4LGiOLOQ14CLuDYi7TU1hox39vD+pLjKPLtod
r8Afo4xq5vJFgnifbOQ1FEtAwzTPNTykQJpVKy5WBYfvsi4pnnn+KTZZnzKHscGY
7+AGEcavjexF3InvKRmaRS2JrqaIM4qnSuXdTndOgBxtOsV1PM2x4DNi/3SWgChe
9awOAJW1F+ZVqwyqyItk5Hjigtq9BpTJjXkSzIp3n2bmMV9KCP1oJEflf4fTBidc
49TtLIy5w4j2p3cHFNgOIl1dxyeO6GlJKi8Ub20wgkIcbfylrOlV2co63AE1K8RR
uaN76I37qfZpcGPUnlqLxw==
`protect END_PROTECTED
