`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SEolkmmsEBSU5k417OYDipNz+aV7O9MwkJhi6oxgrK7lYXrf17ysOMgCApBwed5l
3Bz0u8YQeMwrwOjV39UiAZk2lndmLuA2hJU7ZlAfLPr0lRXU38pqiNVsrA1mI+KT
bHhi4xIlvea5xp9GBvwOVHObTXK/lkCpwyzFk3k60NzpsjV3tZSW2kXFuUjZA7Vk
S0lsBKRAI8WcqOzF5d1sBf/uO0hJ+xDTCy4wpPWplEHo9bSuCToFHaWBaX5JruYg
mwe2GJalPU0zphui5wR4bb1xS4XQDU33fpP5fD296muCySMzr6x2ceMv14A/rkMU
fhTS2w0CpRBnqtHEXVZ0+OHsYuc3lMkzduqXqronSnfgoopDhk7NpCUa2nevavFD
XhcHxZHKuFDBiBv83S0q7+HJGcVmA7ZcSnDkZvYnJJQ8BQMl4BlXLMb0XiR9zyna
cLeCLnwVNirZJ8fN/BFJPA3Ns4qscm3xDHlEmHFAH68l29luFRC6oTsH3/9btqxx
JqJXYxUu+tXdZtHkQEaAeBp4xhXHz3bVdbaDguzccpLgiT0UYGXcYckwz4+wh6qN
U0+eCgeRR7GkkUL5YUZK0Mo/hxbhkx1ZA41z+uRjMxqqFaky+A5I2qBlG6YDPbp4
Rc7K3KW4EbYQ3uUzZdLeoqVYJL+RRM5T8JaPQLH93uxdCcelqIF85KsQg7IkQhZM
iEv8ySq6x8NL1MpOlvjOdo55rjTOfeCcZKMB4MGphMP9d1nkByMIyb9HQp34xUuZ
sSs1khI3IzpzVE/QV5MSklv2OqYE16G9YCsgkL2rSm+yxNnmPverlT+y0w6OuEhr
iB3RR6cq4zdYxSBRcXQinmvdYrJNQ9x3hGq7KhxCl/Mq59aKOahSIpb9ST8BC/WF
tht75MmYDnl1/2BnaJxoVuqzGYtFk7L+cwh49u2fQC0dMcbRMpoO80rC8PwEqh/o
1sTcZ+4Z/kRvfsRXbbDTBmPymTRz4Y82ZvKIYXmjAiteM+JmeGLDcJWM4Rom6ScI
60XNEoxm7XzwRe5dXc/w7laay+8nSGIanneBvGka0tiBVpFr3Ynvf01BkTyJE0iT
kc3TxBQGO6bVpwYMqCxh7TpvADVZUj/EETgyIsXcFPK9+AbeJL21O0xqsQFGCixx
zaiFiXJgvR1PtFZFZVq7Zq3kBiZbmMbC9VZXRRENWdKg3dy3J0aY9hTMmPaOIVrT
GYdtBWk8KPI1kGktIKtxM6wyfOiSVZC5o5cS6iisuhg3vWTQUgLlTkn6Tarp11Nc
sgE0RfjiXizuiRuH2M9zztAnTPrm+uNP76tg7Z/K1c6o5ZmrMZOW3gHKeOGJlwoW
Y7zOSvWzXsqCdpGLd6veGtkbhdknx/G/6yoO/6ttz22et1nL1Lm98FIlHfwqW86w
gJfC7fxcBz30jAOqmcwYqwv/MQbK7P5phJIzklDePwHQwyLuR2HlvyZzA4sy0qcm
RwXPchyGBMaKJha3rU4Uibji7anb5LkIz7Pdfe4+7zfz4e5I6zQxCvVGOedJ1L0p
ZiOEh0lHoxnVlvHpw1f/+BGqHMPVYjKcgHeqfzwYlaFluMqCsDIuYsFv1vv9d76m
9URO++/q2v0w9lRdV4ce0M/h6+1txF9GIcMnnl9SQl74Rj50XP8NxR48xIEhX/It
1S2UKum0ipxqy1juhmicnZnjkE760J5cYLMCxH683Wgqf6F3fIPcvPFMoZjxM1ac
zctrG+EBBbhiKVV+ePd8e+pkxH3rIDH5wKQ2fTr9Boba3VU8YPFtfsxxJibwXVAZ
r5Hvu1iMXQ6rU2UWRl6aEZs4+mfO9lgqtDCwk1Id6cV35E0Bcfkwku08Q2A6ObmA
G4EGrgam0z/isW5Phmr3I5mc+3jdiSDKm7MbqN6sWD8FCrVZCznAmPZfvZWlzoS9
0vKaEtgpPfvmqJkAQL92I/5eVab1PvbKgHMJAAkNX9E=
`protect END_PROTECTED
