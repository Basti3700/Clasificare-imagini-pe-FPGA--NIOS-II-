`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3HK3/Zpf4UMXFsSOhwRuEX1cmalRPvi9uMk6aMJ34My3UOBoMzbSBnt1Z6hUP4rE
mqXGGePUsN2GnbC2pPKcMykpFFXWro7a8KI0Yj0SXBeZy8nJJudlm/N6StXdjVlj
ilVZdTFPQdgd9ZgPEPqwTYjm4h2ALYfutpPs+N5hwHXJOa/ZczNHVsjFqpv7OGiU
geG+k9mZYXXUPQF28QwfgCHAYAcP0OwmT2JJEGxARft0vmuQ1eBay81Q3I4AAcne
wV3R4M9zm92zuSs5A/CIpiVq5wMcZwHYnHwoALduz7KjVxaYeBsn04E7TTo/vXJ8
uzqIV2HYlyCZHsynHS0wKomJV9fz3i/Vf3VEBWtj2/cReNDvY7ge2+3zTpdLkNup
MuVtYcvE6H8Tok10X/yb/TjQcGjddH5kXCS2sNWDdOi68hJwMihKBoup6ITmKhlc
tbVN/5on8RMWl6vm+sfC5tDKjd76mL91Rmurf9XZrTPx3EfetncCdzZ0k+U2fEXl
vR+Vt/j5wMtBfBKa/HdNwPUUVIVPR5xc8Id6xfLsw3wuzVdF9v5BVFOQq392BKue
mkrbEWSWmNbKE/VhUAZt0Q==
`protect END_PROTECTED
