`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgKnTye6ADZBQqTmLBB39XBSLbP0XM0TKRQIcNOwMeSoZjCina0qHuNCnnuUsv2G
VMoQKZb5wxFKU75+teh7/WlozyPVINiUCm39/C1NZsiDDgr8TBqwPlQ/8pWk5dnr
Gj9+n56Riz7DxjE3gRJra1uuCzlMPkja3i2qGpIuYvSgQmVRRXZp3Qi190IWqCn7
R3Je34E8uMf0/pIkMgGhrUmr0ub1u206q9aPeLj0NJKl5iLmnZ5HL4ZpxADRvqQ3
G5HtI2Mz0YgqEozJAG+m9YZ0vcEFUVKMqzDZT6GQoGOJaApzan+d8j0yfEHvcBdu
3br/vKoSlzvx7DLVdeobyliQuKXJazBOfYsiMmWRFu7sBKjZHGi5Ra5EcIFr78LZ
QzdZZZFRCJH7dNtANkUsybAlknigt0L4nUh9yIJ4edpBLqPsZL5iVm5EOyfYmaOP
oZRNSUAqkxLsWu4ibGQTQd+NHyA5Q9dtiBvbB/LJePo=
`protect END_PROTECTED
