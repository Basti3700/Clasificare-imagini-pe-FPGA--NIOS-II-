`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3MR1sohDu8kDQyt+7aJctifhcRUt+ZFJrDvBLiqOnK6xx9pDFguiN/0i6kHv4ya
i6b05BED0TXtkh8mpJ5VaHtoUWBR2z+yOG8I1t+kAjOrIx0ar+b+ADeYBY0YZreX
yHPDbXMbm2j8XgLCs+NnFaVDelergY1f0YAZnOhLt5FKquqLCcULSbgxtUMWAyG8
xgwTE56029s6VW1/6Ckb8++ZInvBOMWZRMhuomb1ue473zKgybImNtSZNz4KoedD
`protect END_PROTECTED
