`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A71V2q+rd2YU/jYBDJZLaR7emAw+KS+ocVpoekr4A1RaiQKBahoCl4NB/FYXcclm
jLeputM1yqboVPEpW08LoMLQIyXvnVdGj9LtcInC+NHJ3EzTcHatRWMu93eaqGbu
eBo6Ua18/YjY30+PPpdZKAxB9a/QgtTbGbwCB+CpHGtTBkN17tvX/xhKMZ8KLAqD
yTMqtPQA/zs3SSvkWIPLtOJTIzWdwC+Izq0DWmUhUnv7giWNkXJcZK5pBY/1GNO0
qI8Wp27eKYc0CEPPjx0GVPLrnZXZnkcd+X7Z2Dzeaod06Ogk43cZl1tY+uYLRNHs
ulHUO9qRKtWbBa9QNq6xMyg04kfFfl9sdnh/eAPwIJfvwWZbasKhi1s/b2HiePck
wMSJvuTmkAkcBL2taN4mbWLxtHPSIEDSOOBxxd9nwnunuHmI+lOXj4nQecHy8gBg
zvWvRjmujkv88CEN4zLGMWSVxBg1LZDP4CqDFKOZ6hz8MZV+W09N/Iy79+bdy3EN
L+9kB+x0N+M9WY5xjmcdFyFKOm2oOI0a4I2aye10cCZYuuZMfMAUBwTavdhMjPnz
3q6ceP8r1/Lu0T/eBzlSgBVl5ctZDB+h4KjHrG1Y6odXrVvpQkN01GO0AYI+P/7i
XbS3Yn0jM89sXH0wp3zhuOniV+jpVsq7UDyXq+grjNgJCnuoj0K7VeaBzbhk/aDK
S/pyUILNa9qYWVlyfYqV1uFUQrGQY6UUPAl2eVQvyrqeQeJqhJ5jNnRYhd5+2Fcu
A0WpIKBiklX11ipscFpzhl6rAPzUcCVedQBkxBKtgFBvOkcpaicf+lBGWdsNe+a4
1VRNAgzoOZ+EGiWA4ArHeg8CqW46OoWDLnP33iL/Jda2EwWtcR0GFYWZyUZ6wy1A
lUts5F0Np/Ms/JAeYXqybNnsWOMJo+oz5FR0WWHGlm8le9muJs9gS6294CEDkFDk
GHuq5helthiZlEupWqEEsqHDryxeM+zKRYNCj//Sgz6jNfgu6PEi6mBi3WPhtPzz
zlIlVYfF8/WHZbxqhU8oflufyDxKPM1VWK1E7AwOx71kNR1nsq+NwYC2PeJQzlp9
3G/waYg9Kj3KIwGGo6Px4nstIfL7RXb8cAs9NlmHp2YzNTRFFzDRFKEyd7CIWm6h
hyQm5QRA1IJMXsQ1bKiNgBlMFge6CIcCDl4ExQ4fsTkUDSAHo1HOimfl1v22iPCp
/bx+vCe2NEhCNuqaXQTmJWVIGwnKAR8qCLvMTAidxtEXfBX0BxLjKLs+1qMkA6Ip
6svWk46QUVm5n+8lm9YkkXAfpsnSF932j61FIeeWFcQdXop5IUFufVZbM51RF46g
Mt36z9Zb+ONQZcUJZXPk/Sqej9akW/2+aJhkisw4gcYtfWG2QEC1+kZ7Ti2G4BI8
JMkB+3/gVQaPYdOuoXDxH9BJnfjnlORevNpOgn2SyxZaudz/bVivyZufe8pIBRZ7
QWGAbMbNjTA7h4ogpXfBgC7P6XowFCmdYi5a4fqTzNzKWlW7gZ+7pY3RUDucA+Nz
v+lzk2OSC/TSVHr15/i9Dv+kLy/r/d/QGmk3iA+mMmitmfWOa7oPVYys1F6T26Kv
VlEcZBLPukPWulbFB78WBT4uNSNfE3jawjCsaJ4jciGUUknIarWjF2ZMpXVgSgW0
rf77dZxa6YDD9wgiDe467G9OR/IBVlGloSQbd03X8JMUtz4x8fSSJVHn71Fpofym
faH/BbiJmALcvtdGE1IfsXZV6VCGXDw8TD7xd/T89b+oVsspWtyTPBXvf5mgrUl6
LoiKSmgzfje/wEjGIaQ5yR0FWNPPPki+drPySudPbWb+ZOiQFCdkIMqVRMKnpcvL
6qTetQqx0Xfj4s6qO+z4Ap6H1uSxKV1PsreNxRagrm6S96he2ft2OOvZWSJnhJXs
3f2uHgCx8UI8U2uJknVgGtCfWx0iis72dZ3VpQWt6Z33SXtisLCkFyfkJDcAIHET
yS5PuFVNSZyCcZHdDkjI/+wfWijxyhWWZyOoE3OZBr9OKafv6Zr8Ejq2MBGNvKB1
aeOLKJsf2rQ3E5Y1vgrfWzW38eePyOhz9mmfMyhkA15w83rR/MLJceC6s8JVgnOC
iQT57QhE+A1z6Hk5ltOUMDYJrd6X2TXIu4xgMWEV4RidmooensDKRxGit8SmZ7wF
pUOFEFlvlfaq4LysINxO8QKU/nulXjBS9crZ1thuZ5EyKoLPi+ssS+NcVo+ucTDk
YhuHT5AI9IdwZeXFdQmiZd/fxiCmjbCm1ie0rqCHTn6Vbquq2TODUycu/ncCbuIJ
+IUFMu41lgjevUcQwmhw+h//Nh9W3esje/qlsnypXLfZmu43MIx4W/lPZ1rWVUwL
0+TuQ0Oxd1U1UzTN+V2yPtTqmJffy3vm/fYh2yf9YmPOvW/GHJIwvowP6sGaaerI
9wxhz13OQOu0rZOyZbgoyNgWkqUyEYIFD2W3NTFLcVUoPx+IN+EpIW56vTkzNo8N
Ncz3ggtChzOE3nWHzWHVlU3r10XrpRa/x7ogefI/rKu8ASVCZPZ3b0mt55p1IE+D
8pFVQXp9B2ZNZZW31pqyd+DjZ1tjzNFdpHFPamUEEzYomCLtKffx/fo/8E5BQmew
vXbhnf9ocB9k0WV4iKoHOacU7rgmMK1umN84h2D76SWtN93KttZk3it6VQMb3gPO
uTZ8VQj6qJAfbf0YjVAmUjvoD4W+1TekX29VYHTiorDoHdtQ7upCTLq6X22akc1U
AWGb+APT73hD3b/zsoedowOGoMU9l6HdlEd1hUZzKpdCKL4/s5CFJLC7rxJN9hKr
cSNXM22jz0scEhV0Yr1B5uXE7jJWXT0wwGWS04hNJWPvGA3M8A39uhDTLZ1Jah7n
dZ026MexhPT3IMIsPjkOfNeTE8Y7YtjxZI0380V6STz5S4Gz3OH5iYDXyW85vJDd
3TA0nguLTIMynz7Y0eJBIp0CBpKGTL0fWv+X796BpuA/B4JfqRK4ddAAu/BxYIPz
eyLrjsYoaTvKpVJuF3ahELNF6DUquSbOaOz9wH6OcUp+QdkKucI3HJl1xc/VS2L2
S6IzhMj7MO65dsL6gs8E6/ZiwRujDYu8001XaqSMRQt6xEz0zrU2Aq/wG3/eSXvq
`protect END_PROTECTED
