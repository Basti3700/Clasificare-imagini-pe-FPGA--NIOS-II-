`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
er2dhWElVnpzHuY7qvhw8WkLQAgB74DH9CcfQxDNT78cAHRPU/0qoK8P5679TrH8
XNoYNYhp/i3GuzCMByUKmyCiJafSdgftAjQbjREmMBCf6GZ+DPHuaXH7nEqmDdDN
t7J8K1soAX0PTn8shpadznVHUTBrR6ZBxVRg77T+mgOkR67Vztiv3n9HYFPxJgP+
z87IWFkpiVhym/KuaOy3MunwxcGGmlPWHU6v1WqAgAVRgQCOEYIzkJple63E59mZ
CbwAlqleuW7cz2wa2wC7amvkySDuNGknYKStEY8atHuMrUKtNu2MkVP/KDopQL3n
3N+UJfR2BsHeeUu7F9h+8TROmdBJxgDXK8P5B+i7yhqBcgFRWD0Mybp0qxJ8hVD6
LLTe0wM0Wr6xfegsqVmR0YmjkOe8a17FVGkikfwFnaJqKme4TNJpEBLKGLxoVo3d
UBicU5j8jPvoBo2b1p/LqXR9aaMwPl3pz+BplaOS3h/tBOR1lZGY1dnqKDvbTTwm
bZOVH4nB55DGNt/sTzZPX1RIfxos5Mv4RIjeWVGzGfSEOEJJ4dtkTbksOLEw/mBw
8FarPofmiGcyMmYEikCILa2B5+HhQJVKZBpoGVdFGiPISG4rykPTklIRvGixVKTY
iGJoiEDkkAsjkZvWGRuzVlwa8qaOHGSaJvQwQ7L0Bq1I56IQqswWSXAFXl8BYS4K
7fO3NojM1jGazALLlhszHaXTvnI8weahDZE4Ls7xda5NwvHzqfSu91LhdYUlWkxu
y9iqLRhcmZ1FGhBsg+2ItwMiKJDOWrpSb/4RtGkFcxTNT9Rp2Cp11muZL5eoOuRy
OcPL7vIron7IJHw0pV6DYnuOltGqLKIjGW5UJQnUTnyjfuboLWPFsyNePd206Dyl
oDpFOrziiAl5g0agnk5XmBH6tKuqXffieBK/d7RmBzu71Q/oTA6wChB3wPz/dHfb
lo+pgMuhY31Ui4GSOcTWDPK046CxJ+Tpdc/VdTybJHG7stuMGGLv23ci+YwDbkTp
+Lzu27MrF6MDBrAx/6QGMglWi5cgpvJS46vXsZcGqhMYwb/KvuTAAVpEsF1dD+Z1
pC7971aLwDYDzIHkPlWNQiCfV8pXoPMLg0d7qjnnxKcRiNh1e9PvFShg331NQt0d
db+VlRjRECzmOBrMdoMX3BwJ9O/0Ry0wIZV9N29CStwUl/WXsC0P+79Bqj4UrURy
/BZBhmvdVivceMsW8PjsfUdCLWHDvqWIRszTjSENio6ryxaCA5CTJoSEAxnTIJfA
399dr9ahSoozF9EycfC113OsiM83crtAwQqIuGuGIdS8vOuGmWe7MpDcqWkrJdab
dsiuVePalNNfDocmtqP1hI2fA329NOCFzi+d6XI7093+BswX4spaaJ66hsbG1tda
8a52Izh+e/LY83RisSNTJU/fRQ4OqrSjsVo14hoYdRicdXtolzQ1iwrqufyK2frq
5PofDn/MCZflU2l8oexFC7Y+3+7slmJLZg0qyvgufsmzqhLhypeNsTjX3aFhoU2A
YRZnQ/qzTlcifS+4B0TzVq4196/oA/Yyb0K+zG1RkCbthyj0PuwYwdi8XW22xs/u
jUc/sTnTA/umyxWxU+RCp3IKMBLf6tIvFhuIBPLtXcDkwzatfAQSBKTKQPtrKxn0
uVF2OXNlzbfSX80WucHw02L18zIe4pypdgIP22iQXWypvvNVYLTFbfYqVOs4c//q
6ab7+U/FAnxfb1eiW8ihHBhOiF4Y7I6dEZNC05O6b8YcBVqmMh3dhTplvARGNdCE
REUqEJd1MMkkLHnk2W8/fRZxc0rrS//oxL5u2yakRQvWqY0WlEKMTgxLz0sY5mMv
LE9X7Df3zDYzTw5tWV9WUEdQkzG9dFIaGMpI16M+jurkkv9SZFWAx1ox2xGE1MrK
qzoBm2skFxIpU+8JtI3+hWdzspdGxX5gibftTbhUGsI2txcBin2lRCDneroE6MuN
zzc7bMX/EVMN+Kxu/ccxDokn4DRhouWIY09dTFvbJkv6iodZ2gIqDD2EWxu7kVj/
WP8HY78jSg39BIovVPCath0aaMKBfY3tsJNLapBthzmGnmL6CLkXnnsgYxcGh0wQ
UE9XmdPj+JsK1H4h+ADnANAx1g8UVYLEagyTv7KIFVkCcqCMHt8WStGX6DUxD4hI
w/T87EyBWiqnkZmRGUbYzHhCv0l1r5bELGK+yBjKEMK6VO7Aw3Tl196+W+gWsp16
E8SZS3+AfdNv68MnDJ2iOsSSwLbBfrIHCmoNceAFe0ojqmmLDcpWBc/1ogDghIO8
9rTGVQbHH8ioxGkT/ZVojzEbpQHFoINQAfBHhxYOraF8u9S2IaJl4WT4KpXuhlYL
79o8fsyCJFrwVZk3xqM2MfsAs9hwarDFpvEdnUD5tVyQyfIpAtpzjwXPNNJFQELR
j/pJDONYWbVYadabmBONWpb062IpUGqrHgsc3sIvP2seGupWYzbyXG0LJPQvdjjp
8kp1wunbKDu4lFOpbtFTiJhh8yMvZJQiBYHIxsB/n92aO1AYmG9SVs73nVonXNGr
/wTJd1LvqSki9z0RaDVlc/7eD6YkmfgeK6HnuCDrBWLnTqU4XzAUBFac/OLlUDMN
QrN7ekkalU0j2D4e+TbNShAbxqsYSFUIBtMjqa2to/888VIheLmdgg1PHMLkefgR
R4TSWfvo2lqZ69ISAZew0v0xFm4sm0q5H1TzThp+xKUqL4i7Tm2hufE8o2smKXw8
9xhxOWEGQrylLEyFheywOjjNa6weMzjKZnQpSfLCT3SrwO22/kbx4k7Tu3Avda1j
hYkq9TkF+NdVT4y4ObPkvEjSRrdQvfu2leSvyNDGJL+BEPwQNeDpmZAY17HLSpqf
8MmhZWpwyDHhAkFEJ0VcpeC6YHvsFKXcOegCujqciCnx9FGaBoHZp3DATZRcCi9p
Kc3qaNNN5PYRlj366pqY9q2xfVOeGscKzy4xg8pkAJkAQsQSwW3aftPRh8p2iME9
uItfpkf7MJ+tFloG3aw78SAUgYw/m7PEADy+Dt02pHxjeig9uUl/SY9YguLkjyin
8MBP9pA8QdvSCKozzt8zbmGyDi7HzRFX8/5FKiZE4TXXHUj91OR5XecsCp6Ap8od
3mqwc+n+27GwYvbP3E2pXVHw2v/vajVg4IfdftonRo+GZ8+zHTZf5J6tvAtpVmwL
VqKRrpTOJq7mmRbkn/pBa/5i5WKPAxIflJuzlgpJtMDcON6fSGDvmdHAZZiX/Pwd
Cst3ijqgane1E3XnAk0LJ0ihwrbAqBjvQnFbzRWfJZYNNMStIxV4rmdQ5O9XC7y2
2CHE/mgjdgswmTla/66hBeXeRP9J2KdKbubkkg3AP0U4NXEYiXZvI5tsGLs+VEps
9t/90Kh2o6GG2JgxyI3K9mRG6whfKBXp5TlE4LEMT67LSQlDnN464OXua3R9zt7u
s4H1Mjs0BunVSxJgDLe++HTSdKByPMzLaJHPggkU06wsfgI9QtBiDNoQ1uw8TKWx
D82k3yxxTzmF+DHpFYug/4q2mt2ulFM43TAx9U82KOhgtG6kAcQhRA+gsO2J+9Z2
U7Dt9CW5kjVScDlCAMNGNzs8zjQqK8NXGFiKCMr06Wp817xWxG9D+nlPUlzPxP0f
Ot9tLOJHyCvXWN+PB3kUbja4AVq0LxelH9qTx6orNzjqefhPTWzFpnft14jMwqVA
qm6aWsoabtIZviTb73IR5QCsqxV2RkaWa1pO4egLZNrHMn6AfhYIWJObwsWTKseY
qxoRPPgY5uZJdPOefnRIKYwD4pTl1xOvZQVdunnbUk7/TYzzFg+85kqxm4FONNCI
XV5F90La7ouTtibadTy7AazlD6bg+mrUuc+z8cvwTztElQMim8kMzlNpaXqSlXIb
dD92WgSHMQ3ACGzFFTgMtl2KpwK5ZgvO0A/3Dl1p81yBpvYEGyuRC/hmQEhqaevv
kTfpwMEHIxPzcAs8FZ2nq/5f4un1u6McJDIH9SomRgw8xBQ0TjzOSOfhOyEp+b8L
Axsjijx0wH2jTjG6gIWLll3P/xu+qtHuHW9Vdx06MG4lkS7kdlEf0GWiJqkH0Qhb
HPeSlbWddB9+iR/uCBnZoukY0JJZTDdZgsSwED3mBu6lFWTEqVDAE6xQS2kkJYEn
a4Y102crKlRRKzRzWeDp0Y2zNEcZR48xOFeiltgYBf3w2TLFA4BYo6R+5iQlYnRu
e25nbKIq/EmC2BcdfwiyXGomkRrtJ7lXONy8VVf+93a26YHeDjVaT/3yFHO4hqzy
aB8cOIl3aEteS7kkMxaCaNIv8sQDSnM0/j5u+2KVMlWACiKVCJPjlB+hQfS00v20
cRtnynOQOnm5VACR1F1DmDUceAA0bZce/vVSVy4kZFj661ccY0RRut49ielO31HJ
`protect END_PROTECTED
