`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
merMspGcpkzxcNqYahgk46MzntvPrXG7dD9BCBSkMSXMAqzhwzDDVPQh+AIMwJD9
rmJfdlD/dLFcMcY8frUY/rlFB5MrJHW0utpJizJB+L22LCqVXKOjf8cjpg624y7d
Rn5OL18LbzO8ek6zwgV+1c0xmgRmVV2Zec6QIsOlS1PmX1Pia9uyWJ6f066UpSqS
BmeKwlDWononLWmfaKQAP74D3kZBxC296X/+W/mWyMfIPnOt/uu33HwSTNhY6Tro
`protect END_PROTECTED
