`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KLMvtm8r+IpRg+ySYTh+y3yCl4Og+rYajVDjArZeOxB+/9WzuGKlYiH5InLilzg
2VS6IWD8aMJ5vZa0W1BhvZugArISqeLSsxgvMZKIeezf9zRL0JSkHKBfTXFr/NQP
Ip8cgbG/wbnokaZ0XzYXM3L7/5Ra3W1rRYU+sPYXKZLhBrictnEV4g3odvLXmXkb
U+gKdHbj/ADwIfICXanpLYetFR9PVYRTEU7CFYCV3W/DSY83mwgqKH6nWHbwcV2/
TBvGHrbdaQk9uQXmGuQbefIdlCji89fA/qwQSEauTIuXYriTX6l9vJ+sBsfeSu0u
Zin+Kye61d/+CH51LiaPdxMW18h8ONyKgrbC/zTJ9MfdfDYbRptlNZ+hsBaW7gwP
`protect END_PROTECTED
