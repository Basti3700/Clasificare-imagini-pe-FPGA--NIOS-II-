`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xiw8GF58IEDrrQM4TOXgGlmIg5+iEVFKv/tdOiJkclgTomSCGrQKiMEt3zAXhobS
brjptearOl+LQkINaLtwwR5ToFq+7i9zx7VnsWXbpr2/0H+7tXPK457ugwjkT99S
1PDrT0iK0pEONRbYywQSlYba2PpdYj5JKU8G/QbsbxwhAySsWN+19ArPzevfPIbN
BQmQuvHugxAuyuB+SsEW3+0Q8+WSenFBpRccFUh7tHaRtzcrjqzbevo9OrTl+mcS
5sUw56Y1LJRYnTDR/ixVFrvJGPC5TdTCsSjObuRdruxcxL4LbVCpJvgJcguxSUVD
TrsQlloiZ++MJWB4LzgIKB+sPJWy7jIYZJmMKnoH8mnysDSVdcmLTuaUH0NsXJyU
KADaHoTgyl8M19TFcVeL9ub8cqq6td+kD1IHz0ABzp1gyKvToPczpfMQI76PQ4Aj
JDBDo1zgt3SPSMVyWrNR2ooFs7SnYPnt17QAI9us7G1FGV9Njk0Q4V/qNN8VXgek
p7voAyHorwQICOVgIkQ7hr6TmUvHxup4m6AXLnHwUd3WchAXPd6doVSRe+YAZgFf
tQEIyXgl46ep9SKA92seMiOyT1hTOTLU0bGVwPbKXMRAakKFgZrDE8+JWY3t8OBa
T9FeTzlAwrOhdy0DTQyrxSjTGE0fxl7XqCaDU7HxC14E8coSs1cOV401VqRS5rxq
3syXWf+A9l9iXJe1LOIZvWyQwlOOz3BMqhIVlMC8lkvLqqb6WXWL7EkUJBjgR3CM
Ouux4ARuP56GcBk4w5K+D/wgRm9f04hdLjH7BSmsXYEuPLxZyI3YQvURdmaGGpbm
v6SfcG8r3ZUHN8Bjp4/UegmSw7jQHJmkbZkCmxnWfak4G1H/pZoYYh7ahwBvCZXI
kKBrIWtRd3/jnY+dLN3c9pWm8220h8ISqIXeGNTkwdXuKW1GqWTaY6/qnvF0RbSa
EnlKIUQmySKrCWchg7HgRxh5ITfXGW8d1pq+ZdaFGJ/ZGrOL9d/xT0o+VwnJNo5R
QUcBzUKDm7FtmU4kXOKqXyeDvD93GhkJEF01OQEJijx37Ffa0BRegAtEapPek8xa
8bSRDEeAWeB+sj30a+adHEb2QRaprYO9jRF3VOVA4jwxDtgN2YcGv0VbIcSa+5QK
7ezz0Qz1opuoII9BQOQMQ3TSMh+ovTDYXHc5ZwDbTIeaUE8jQE4mvAVxcbTPSzOm
TZ/lz6uUJa/XnSijXlakuR4Hn5ubekzqsOYUDfz8MsQzgNRVsHcnYi7oPcPGdREH
UkbpWrut4h/sM3VLEIN7PtuctzOiZL5NZ1FOe0vdGHMMDJi4soGCHpk6CPU6e1/P
6/+3jlkXmK3GqS5aJWMrC6FjHuDfGyhKSi3j7BkMDpzP83QTswF9NnHo5v47luRc
u6Ta30gnV1J5M+81s1hsqcADObexUfEhqvKDqq458N4hDhTz94dQJixj7UkP2HrC
FD+C7Vd8ZtpOIfFxvrkEpg==
`protect END_PROTECTED
