`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8mD4AtvnGwlw8Xgygbks//JThZa5orJHplndWlHnKEYJPUIbJIR8V72zwCxKOEz
QuG/lc/9qNR8edwokeD47FQ36pjYSYas8utX44BRtkkGVBIYnj+JwmRYwIzq9Hnp
YXr2afircZfZ1hAFt9+Eltnhs9s4fP7qWkjAZwixOsQ0rXhxwzgAHrW4qhDfeqTg
xe1byVPnXKjvH4Djm+6w/f58FSsgywDqbqWsBhWdcTNQUanJ+vpEHSpDYh+qi4Jc
D2JxlD83t7O9g2Q9pJXgiGoP8bZQXs+qexePCJEP07QurVTaDyt9RgV+skyw0QER
Bc0haDvRnlBJcBOT2LXanwZYiA2/m12Sf3xX68waP2EEU7JWI2aufbsXhAGbiPuZ
O/0BJT9igO/0xyDuVRNBHCmWFPnNwwhfbA4Y4HSp74TKeijeonbHPvCdr5+Rzz2s
XeVJD1jAeSs5uhRlx+2X4w4yaBVzjyE3kCZU0E7qOYQOSc3VvkNKpYz0AGqTgOWX
fyurKzzrMjYzuN6X/RkrugMktQcncQKkc2bLW7SVWSWN5ucnMR0VFbQW08j1jwLJ
Fu+7XveMdPjFn3yM31MpU/PMG1fLdwAxHL9CoGVNpXlQmO/jixVrZOoAaZ8jqcKn
EkvORx9fioygpCXb1wpsobBBC1ooluO9suwiDh5hQK12TzibrvXmRsDKrtf++BAp
n9Il012aZdj+Nm+qTfQIVtSj0lDFmStyJOxnXu9JJZVcN1GuM7Hb9f/EnwvPB19J
ZmpiiQmCjeR3U8VA0ZRZIZWq0Cmna/tHaZi/GaKFHJ/mZyrpnAaWBolr3HzD2MHZ
gdE7sQYiYXkXWYsj/hUHYNwwXaQhxD42pNiAZuJPUR4fSU12TZa0PViTmE/Rzj1f
YW9aEuiRZoKinIUKVsFpIju8lV79o0zm+78PocL7RfYMBXSX2ht2ay7tBJ0O15/0
roLmmKGHedWVmD5prsFtC+1I92iYo6mxcRumXWDaejtyTGhdPcxkTWRwRkXhArwK
9/ERM/aHbkoKTKZghxzd1tdcTnyH8RChgJKrGMrUxFHUrADGdC34hFez83CllpCY
7OLbxhrcwKfhFKY2siJUhGvq4m02/an/ptGDGmYxIrpFK1UkHwNNKJ8s+/M8xwDi
kias4RWzNxqy+jUBU55ih7LXBYDarD0mQtG4W6UB/2ap+80F9+/XoKOmrmn4XfvU
iLdzrifKBadMTThxNzjsmbpS3yT8x4KAtpXjTHNhglawLkfPNlNa81arwl1cZ3d3
raW3eLu4R92IFCS8FdtOEUICMrcVjQNWfQvaqphHNweOLiiLY5YCADphHQDTolBF
YiDCIcTMTtjDypV91po/ju3Y68p5qWLs5E4NjZ3VWgjie0dSyvl4hZpuyKQur/Uy
sJcBUQ9zASeTmi8+Lyqf8MyilpMGJn/k8p+PCHBvNzo3HFb/y0n5PJdVMzyeNpc0
IxQEaBiy75cP4a8A2vcTZUsb4qCNNHKX98nAGoC137xeXv2mKLB9x6SK6wght8mp
VwHMHgbx1tw2iIKoJ5npE+lXpTmDgEp3X7t4y/k3Xq73VBuMvGEgTFLLQv8mdqog
jsPJXlRbcfmBdVGPBP+sE3KmT9n/wjDaZc2INwA/JWGJbW3mcXPI+p/d9v6GfZnG
wuq2pPdNWYLk3imwI7Qi6LTuzgt4M/BLiZU/qvZUVJYEI9+TyuLPXKXaxNqH6mmY
qsgQdJH48Jfg6hoRYSkdpV0j+KyGfvaNGlCgKFaaBe5+I65XN8UGMOBabiFS4xKe
Zz7VuGyl+vV9nYUBEOdMvDQHa0sbIuZJJBq1qHFck3YMK8BjpNB2lNgH8UxON6TK
r/zPoKchiedJo8PuVSun/LG3youtQJCUFymPWhC45OrX7NJzUoJdbGKvVY8XIukd
FsqBDK2AQD9XwNXkpVzP0lnq1weKCw57KIQ+QmeRl+xZ9qqeRBPiVK8oVWJySkqx
mO/kJFQp5abL9n7O4cju/PDkE5ldwGXQo0QktFotUa0eruSs+LDJoJpDdiP/iNY0
ApgtLnYeU/4TYygU9pyiPA==
`protect END_PROTECTED
