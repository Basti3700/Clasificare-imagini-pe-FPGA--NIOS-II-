`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ianbygMWeXiEf5L1h/p07RMppsX2rbNZ5bcctntZa3poThbMmexx/H9QPRE4/uHU
ZWFbopk+ctGT9z3HMO4+LnUYZHmkO9Md3xOcsTS69A75b6jRdisJ7CXHYoKDLc1h
bDjHPx8UKwMszuunVlov4VHuDTCTC/U2K+NxUc5dcM/fW5ry9dHt+stJByAVA36X
soxxTfhc8qjlwHzB6rk6ol5t0pKauoNquyNsBwR5lZbCvjg9RiYaey7j8Xx495nM
oNUJeo63p7VGBGXk6W1OsIQaJv6VLPkAO5daqTtTUYr4RjdCYwmV8YuI6scCk97W
4+zkYD7agw7gdxS3ZEfrw83m8PHXIpzqLY1JLZAvDuvZcC731H8kSp4b2HT/fT+0
`protect END_PROTECTED
