`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTbhUvJqpYwVE6LIlb4mmBDlTlMXgvw0k/NPMw2oQWa7ZaiMOO/FfdAqpzIfjilp
nzepnNOe8cQumXgERjrjZLRx/RmROImlmBTcv4omWMPpAfs/Viwvb1yYA01jVM1z
DwxkGk2RSctL1pQaDkmXBTYE3XRraNVrm8t8dN6Fu56CXyR9lZS7tran/v9vJKP5
VebafwobxKX5yABnafCLRFLugzFC7qH6/3UPFMpx87kNBiBilsAsV5/nfNpBK2nL
DjZu1GEVcJ9kyY/+xaYM2zhRvACvfs8ibEwHCgFigPmASpJBr3ZsZmSpjV1QxG4t
2cUITmozQnbb4SX9XgiuyfnQXmHqTePiLXCdNMYPxU1mE3LLyxR6mpPksq4W9r9n
+Hxt4aFhswa4NOVOrHR0dkohzFYvmvsvUmPVGwe8xR/BvbrE7zzxuHp4R0Cf8AgL
ZotFYSo1IvXpwtFr8ekcyeSEJTJ3kyPq7f3XVS2RZSmo3C/m56yo5v6EsCQD2L9u
MoSl/TF4JqoTd80t1ssVqaRzDKXDstL11AIqodcjv4l0SvAo7rVbM7ENAtG2DgUN
bNyBsH2KsvHawZUUOT4ypQ==
`protect END_PROTECTED
