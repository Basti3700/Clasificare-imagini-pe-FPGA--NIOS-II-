`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkNppdxPAU+lFdIeyN0sbSSxO3P8Ns3/oLAKSv/YfOMCOHvU16Dv8SzFzCCKYVLU
QWxq3bInwU4BG99BmE5BDoYfotvn6sp6ex+BvPV3q2AYCQyVRx2A+UVWmVuowQ7U
+6NroSjhl09YGATILtA3fOz/znB9eHqsvguUsg8F/eAppVVsKcx3VBXzAM8I6nVl
jK3edSvZyqwbUAof+jF+4Ex4PBpLaA+jjrUCJ54P6Mq1BuX8hP80trrRQMFXIImh
DbFE0QvA57Czk4M8mRo4UkwYnlRQuZFICmMVUzvYW5Q=
`protect END_PROTECTED
