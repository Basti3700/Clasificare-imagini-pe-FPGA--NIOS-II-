`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfU/GMy8fOLH91g3Dp20R/xZiWJGmrZX8antnDD+vDcJA50J5e0sg31Nl7srQhDl
Sckpk33wqXZIQnAveChevXgmgQz8BXpFvQ/QtwT38N2oFsr9JfN7mhWJ9ClOS2Zl
lWBWqeFeP4xb0SHhjN37jD4bIDGOdl7eXMK3EQ1KAcydwnoqjJ230O2xW4ZOvZjl
0ga9rqV4+1X0eqpvVqR2pPK83pfcIM43I/Dbx+VCm27ZsefugfVPvoMa3Y38+HZY
iyRfPrunKWgs1YhsPZlGdVStWS9FrOFktvSSmRXojMEIU+TmGBg5PndUxqjDXg8G
AquwQy4b2uv3aIvihsZIwKp4i999KA01HLuJCfN4m21G0/zX6TrQnwNXLyJtf800
zlGTlMtK1/acnNuelQwjegBQmHU1yvzLGk8WcuGDbQYGYLISnHB+qXGTYGjxGUOq
IL5mUnBG+UxpJmNYoLjRb2OrTw088Hufqk/6exzeX4Qu4KR6mhByUMlN63tYV+wm
uFs8ln9TovFnPnDAK3o4FEwGeXwgGTYgzLEEZ5XFVei03oM0BEZ+bPpmVK0rnHSY
TGzKGD2mBJ7ebPQPdMkpycIQb+a1RX+DVZlEp2pz/xMqapXkd5jQv5adUST2P/1H
JkNPqJZ+VcHTpaI8GdUkT/SYs4o9KyY6q5ljp5HQktw=
`protect END_PROTECTED
