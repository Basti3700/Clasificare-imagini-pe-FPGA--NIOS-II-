`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2KpPUZc4OMzegonHFP/y7ykAbEKdTkEufKJzZhZoNXQGnq6gvoCWflZiybhdQ27Z
+VFgiKlFmDFwgHNibn2LMqFk11/KPwLkyOSG9ukEYs7ysRnE7TY9yZcx8fel51A0
JoYZ4/nrUBc6zzac0tqgXgS28wiY0RkFt+pyHhblt/yJSaxzUsyE5NXJuO4Vkg5X
9Aas22SBUNMk51fXqnoSQu7R4qjxKeURM13sZSpc2Cowg91TIwfDTF5UWfXCHgWd
xyUrpiZaVbRpVkH+X1ZTtnDpTQ0TRObdeJ7SebX9vCmAiUkGQRlBH7R1qdTkVoH8
Vx5q3pTKxXaxG7ajYoZQT0UlaLqGGMHTK+BDgibAgRMPowWzvyRoQqlKuWoLQI0m
2SYLs75GV+9MLZ7vnX/oHBdOhQ82KCP4zXqb6Ns1mbQkKAnY5it1lDv7XnNxfSj4
3V/8nqYU0K7QNhsyXE6eu42faKEvlG+aBPEMRxJN3YSVUVGOOBJDAuIUx9pj+8TV
Kfihozre7zuBpHfX189ptZMF+vYkNhe2tV9w1P9cXNWnasbBephG0LX8fpqhIwGV
X9j4yAIh6MD3kUE8HfWFCa1rph6rsLG17AgRJi0meQpExDIui/sT9w71rpmJDzDE
W0RqVt+2oEWTW3lg7EVGUqmVhviw/kHi8dmMBuWpER6iNCe/JwXZ3Hz7+2M1qKwI
2AhtjmY0ZMVHdtoEyeuLT8PWfMRYDWdM318koLiujAMtnd2jVgZP+t/uFj2skJHP
XFHtEUfwdP4cbEBCuu8+ksO1surojW2tRZ/Hc4lqAYnKqYoBRwAhfs5UZs6IYKs9
vjNPszzFmLxc9tJykILts7jtCN6vw1iqMayyBUwe7TfyJNAbNpYKSEkw2Jmqux+T
f53oz6RVEi8k4Hr7bOWUsBi/ubioaoe5NqVFs7KTB9/242rkeil90AlVNUZwbGMQ
iXGglp2nfi0lXJv7F/5lvYY/r3UJ7IQzLsStoi3d/s6COxyJGHdNAqIJAEmGdMEk
M9ec4ipHICY1PT4RSZnDTM27SOnWhVllq2mxP5Z+ZNYG7fSHgUTofLMjhS+Yc10w
oboWKxdNhFaqLMaoafn48yxSE1HOongunAhq8uat7pVh2xpgox+iWm0GG4OQMjZr
l+mZgiscSGr/lIMKOqOGSyWYw/MuRoS/0i4bM0uh2xWnZYi2zcIarD5ABAwhMnhB
SxEGmk+z6oePDPeRwkNGO/s/mvtKPcSfZOkECtkljtxbubpLIb+3pcgJzVYJDZL4
kHLw8q3I7KZUpj9NiWKrgjUlZqHsl8FSAzgwNFXcDpxjTY8leE0qpc3Wqk1wSKAP
OqDokgoq+qpKCgmYL5dNEVIOg3MLNfqGLmAxszWg7kvARuavkYg5e1FVk7W0Te6y
ozg/25bt+ssLdhzB4Xwv9aeU66sDj3rR61MyXDXE2ZxhawUKQr432hOjN9zjs4aW
HnJcZ9fkmA60Z2eGpfnBQJXuVkHxHZsL4vg3CYdkfT10UWB51maJFzsi7O7+FDKm
eRlsbrG2yHrY+N/kCaecvz9/roUfnGFkEmtx7lD/mXBZoLlIOaxgPtfqGcYZLYY0
4Gp/rnRs0o9CX0NPMM9ePho6VUIpa7X7q0sxjK/0B9EilK5RaZzZvtPSGyd/1JNp
riHbfgeOKr46vKIwojvdxPLkS0czHLS3kaqxIw8/2JkbmTe3lsnHEuiDjctv+IlD
RjM53vIr5kmaJIt7Eu8V5mpH0Z48M9EIjNHGiqX4xCgMCdhVh4zJhf94QuFMN8/l
0yGyfvqu62RoXljrBqbqFydBkmlH2Dkoyg4/Xx8fpTjm1mlSGq/6bYW53Qg9ss48
r+d33d2LjOC3i/YVc0QWcmjzjfBGNqZS359o9UuAcMc3DkVdcf97Sz7GVrsxL5le
hCb+NzK7y3cHNb5xE8aGqf+eeVADLyhm/GbB1tGg7TJzGA9yS50V79XBCTw0oqVi
9/0d5bdId5eIgWDOSwdU2uN/KvNqGCrZYZVaDTljtGFKyLAaTTOW3Ajo99WKPLfx
x4rRsnU7Pxp5YXLrf4urefAAN7YAxcTn6IX3n7Xsx/1a9oBnPF6Ea7acurRFaL0m
kwx7vqtaykL0YGbuBM5Yydxa+4KBxIhRt3luTYGpvfKRRqTk9qqa+s4BIIOiV7C4
giEsykDVtsbuHt7W2f2MVZECnosqhHL4o9To/TMuzhsr31uG14SoGEB7uS9bx8lm
NJjhL+7H/8wGmU8W60PdBtXQAhGSYnulMeaCspZghuGTD2Nphj+pWJ5MWICF5PKD
Nu9Hpg5WAa2zxJDXeChgZCna13PgmWetE9e4xh+tScY=
`protect END_PROTECTED
