`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNsBhy8aFYAP1k7x0kDN3LHTCsm/CSZs8gk3fcXH3MkrUd5vRg5TGvUQ4NbLdwYO
b/hVu22svGXRzNuX8AXTdFtarMVsd3KaVTJgY7ffxFIxC95EWk7rxdwdnvucP8k3
O8Rq+7MNLrednyn1Bmn6elCGrresQ6B8VInRHBJEa17PDL5qs/kh9gCQ4NP/s2l5
3zDWQxL7zq/ggUdREjyYGjV7YIHI/ojIGZfCo9X1idV5RgXdctj5d99YLmr5L9jb
HQXbZ57vHWRZD5U3+D3JQEyMyVbgTBrnQ2lFmwAWyXVxGY9JlPMFbsL0rU0PmaLh
JUjKTARNO+qPf1VzvpDJWcicOUsD7+QGeUdvNK4ct/Xrt1XmEKLVKAcLso9jx/CM
ZGbmDh5GJKK4EI4YwtaabIgVgGxrbEJppaWgMJe55d2dt+I7XsoRLmbVaMTO+ZjV
kseT2iEgKZYYttHwdDOZUC0Z64Lw6K81InaRCIjVDe8cUzsywv6uv1xJ62l4ns1x
uRmrVkoVDIk4rq1M6fBetlkYoT7C04x1U/Z8VgDMAVVwlANnh3hZqHhzJbh/m48W
FMzNKREZ5gRb0mvJerrfY5nZVRcw4pz1pXWnAEaxb8xnfzUUxjEtPl6v6rlwo3NC
VaPsNyfnq8vd9XTYE8LlsV0iWhfMhal/f24O08fi0h8sixW+NOwdL+75PIXcRoWO
KwmcMJrTdxylyCbqwfRij7ZVYzsxl0Uy5cqHeXEP5PjCf7UfqlF/RnY1XVunp/Rm
7A14fDmmxeG/jerWvkDKB2lvZz8UoJdxSoXS34Inwrb7RHWwnNaDu33F+2NTpehC
J6PH6Ci5sR8rrLXN+Kvwn3LhNplBWsivsXN9VSUdO++xZKTkoxK78DHWHRdlPgip
sCpIy8UqHdpjGDx1SuVhpc7jJ925KmOjoyY0qqtzQR6k5O6dLlcTdNGQcNYR3kEN
XY6OrtfhH3kjqkjXN8waGB43FFkbfYYKzKuIkrq3cvI5Ck2mKBFSF6sooferZ4zl
XZ2d+8ubRZ8Gtz+Gx2GvOGylbPTe+ow+yJP26d9pHNk/4YM+R/GPYv0JkhnKdIwE
KmBP14d7l/yBvVhyBV2sRjss879k+n0yWC9GLKRLzQIg440raRoGdTJlWI0S41I4
zNhggNOHereafOyee0xTNVE20Lg0xZ2EltsEVVYjCjzs3di+EskJI5f0gAo3iAjS
ZuAJNcffeDojA8tSoO2DdJiaWqkwyBKdmuwONPeGGI5gS9lhnkAOArLiLY+spKjn
gtcAJPatjOysVp2vO0oyYutT3rTBgWR1U3A7is7cPAZgTHUE9g/8+PRu6/EWcCZQ
LTyjQ746rvamOh1ukb2YR5tl4lUdPCj3crn+Bld8sOtxerMKUlR6IgHQ3lYmvf5D
90yoGkoVcvnkvFLPdgBaNH5xpEge7yfSxqhCg/1T8bK019Wr6e8G4fWRIDnSvWGM
na+XVTuG6x8XwsyD2ZuRj2YQfM2rxmLX1+0luJy1n8vIyX+mUcqmWVtvgobDSWFD
ffyLWG7+w1UPQGafc5IsJNA7D3j+nNkZz48rW1pCVGsTpJwmLCPtInYrB1EtYXXw
W2z+r/wTmrbhDWJVGxxuhfmRShvL1BpVj+oijAnsb5+X2USmR35aZddx9RysaJ/b
de8kwnb3D3tiIDsd4h+saWTJ5v/BOnzDF8a+GgXnyW63YvuplsmyyZKkzEm73La0
98Y6G/wIVm9iahnGSyq5Td/5kJ9vkX+S013JmhD2AbbYzpanbL/JOuM9aljLr5MX
Hi76+gm6rC3vRF+8BcCW8e/w1tRPu3BUHTF7k5EDZtjk1n3oE2u7vxZpTz5SznyA
LyHgO5ODQW88qzDhfKpmWIAXsZnNKKIYpL5QRf2EnGgc8D68L9iNp9drSuPvj4U2
WsHuAO3XXCmU1Ol/FqSGfFrw899YfPybKVU9cCg5V2anVuMmbjdJLAmF44vJbhHV
fGR742KaiedmTa8i8xR4298vuxPExGZSVDXgCQ4HdEHLscTNx+f9ZEL7Xy6ICUva
NCW16JmvCjXy0sdYhNRani59bppistbhxJwpCaGZeHirCznS8jVJP+8fTyqx0Z45
Dcs9EQ2Ybj9B/WBhP5+7Gz7Sdi4UPjjorsfEDA/knEEhYNOOdKLz58BgM9O5qkee
hA2Hw/S7DroOkP5YUV53fcTkzAYQb7L+enYDpoUAyrH+Hh8opD5GP0qTWgCdRPpb
RkKYxVO5aUD7KaKCItf6sJfEnQ62Nz+woiF7D2oJknrJ52/33uSMSxbLfvNe1lnQ
ZgQw8U8vH6jBm0FpeYGhc2EBrSv2GtzxpV994zKpOGzDKbwH5Vj/hCjMAA6HYFqO
pEElqhG8OPoB+PoFXVck+H2imOMmwVbQ1ut36a/62ITR9VSwXpJBcbRKD04Uhzbu
GKe1QTqwW5r9JpNl5kjKraFG5KkuO86MSUQbnSTBI9FCmiSMRSvMFCVQOooHtXZk
rYUAfIMltB640Qv+evaQADu0IVdZwn7u4zrFGB4koYkzyd/bqnheep8SyFuflMZe
7Wa+toh2HYoIEWz+ehrKpEBncVlLPRMgY7iwEGG5kr2trhbreG+DRxcsAY4kB3D9
h5vwDdNqW7yPChhHQoA5MugyTrBMUseS06rxqoIEuFmmUtHnIAeDSvMnnmZFpnuJ
mhgCy5zeDXwqySK2Ko288zyDgzBLOa8yH6RFIKlmPXwf1BGrVDzTTD/2Za9QZiG9
AQRe9InEc5Oq63MoD76OM8IIkg/Ebsi0cbJw37Z9iA7kpppOdJDiSDDIodBww5jc
a6aLD0Ry8bhLMBVJE2W9v42jKjm59WRjQ+rRDVz3z4a+H3gQx9B6u2ctChNVa/rK
CJ/nAfmW6qf4AI+VnKz7nz1c6ipaAqxnMVwYxo3n16QT+JSgt6SrBLyCOFaay5iM
2L2AgQmQidhOll1icYq1GYrQd1TECFH4ig3nheG+pp9ectirtte0YywrAIOXD6JT
6ehCRgKmF8K5nSUJoxuY/15/14mDN8t3AjMKPTzrHImScghp8FqSOG2Q3x3mj5dd
ejz7ytb/42374MUutGOiFzWS1N4DmfTY+WEQYWUYUD3dS23hC1VbcoIVPNl8U+Js
MY9bPJFHWYrwbWafIskcGnIaqJVAHFnZ1ZKWOKhVyRK4f0+A7B6+TMyfHCUDQ95U
Btu+yPVbbagDG9/g1LsahK2A68pLWVcVg5jm0u8GviXeA3e5CBXs3ufgI/LbfhA/
uTlgF3sdGco+xpvA6WvTrK9IiDw5w/ouNsyDNBEk3ZV+J+GQ2077Du8TTs1C6nBm
xm0PEbewcNHvtjYnRAA/Pkzi2tTTIQ9byCQxvtSMOvsLcbAhwK26e3MQenKyY/SN
elDCdwB7JSziCRgPhyc9tySlTT1J9jV0VYYJ7jIPrwSlsJTLCKkV5cjtJsbB73Kz
30v6b+yla5aSU3Mfh7N+O/G1oeGQ0c2e/25GthMULLsn6iiEJTo+cU3B5BwXTstp
LrWLoViYaaXpSjMGH1Pb8M2Vsls26USwdReKgl3SUqewAnVN7cBw1XSqUaBRlRfe
ezQKlZmVAVqUN34CVmsTdKehUDnm378u5CShFTZ7oachrRutM5mam6hq3vUAcR6h
bpGZBL4/SPwnOBmuFHQ8kmxcwokClu6ofWYP+VWa+rxZSN5Eyz8yHaJgHpjrpAux
bNl69g4rmkrDIbV17l4gygq933lCIhSJLn3VNgtTqYtxW8aouCa+cnQ6M3UnTZ70
iZr/DXnJk/ZN0hIkFa1eI5cmObUbyjrr9Hex5mUf8o6dCggb4BnT+rkLmJ5bJ49g
CPzfoQ+YKRVo6v52jOBKMaeVoe0K0ZH1/7LQPmn3HcspKPhzrgkdbpE9k/Wv0WJv
G02Q5zvPhAoVjnD7+NjKXJQsbl0DuG/0OVNb8mSleh3TL3pFchB0K8AB5EBkMeqN
GfaDU6wwTRGBV3RzTPL2gmtoqdmUSkzVxrYUwLknpvkADlApHZ1FtenJ05Kljfmd
qRgOOiAGGvh+csQCOTzAOif+TelAjKnHiu8jHG3H7EXLWSSrxsqlytR1zBM0XnaZ
0htcDowuIzL7Jf3lk6nWvdu5isMm7CCTTqLjzXV66o0Coy8JNhUhJ9h0nWGaMaA3
tbNOjpPFyw9ErdaQKMV98iOmOIAPie1UOoMc3uuRpP8nix4TtQepD+84WL0NDOks
P0e9bN+l6l4JJeZDbDLxvE9Tuq2NDYPM1JEBsvJx37E4f76RQUhTbYT9HL0CJ4P4
xhEqr+Os6JhkpFHhE5Sd3CGIQ28blh4p/0JTFv3Jc9LAmKV1N2V0xDKBx5rLZ/zZ
apOFBliS9oHr9/WKa9KbKYiEQocHqa1iBXS4UKf30Id37h2BlIJaIIHA/kIacn3M
RWJdSQxNz/N5NLL8+BIDfL6aNeiCWKYiysGT6Y4PtPyJzstCHWImQWRB7eVGgNoX
bcp4alji2eknq7i7AqvMOVGQpZ/dfWyySDPlCkfpq3AkNXeVWDo91V+sHsLIoKTy
HiET58eyFhJ4+Lg4VQIJ1U5dwXYbIymsK1M2WKZOkOCYx3K3Mv1zf21VH4sYVQGa
pq0Y0SZh09rGGT/xubL0OYIJ+YiON1Wm7JN3kNY1ZDi3WeqQqU+Syg50HEAqrqH7
1cCWc0y1fLfJqBpCyflKYQy9TYuJxuFqFF8W2ragmo5DnFmiujC9Bu5IypCh+UPu
JsoYskTWno95ERXJDEWij0Si4qL+OFC9q+y3Wj070VZvc/KncIlVOQeFG4ky9J/g
dsyOFf7cqNqA8VdQzJx5ySn6yTdcydlpQe/Ly3fw/tbro6C8Jb2jdEK7eKnhSkkL
1cv/TS4O5HEIMm4zw43zTSaV+BdazkL75zuQPYI5j2OorrWmc53av5cBFtWpK8ER
RwVGqmTwwQkRQvvD33IqpWZEjF0ot44PpGm2CUeucbboBStrvObK6K7I5jmR2rzM
rttoeq5oVE94hocCweq9St3BeujwbGyouJBYeS2LU060PveI4FFgl1B6N00FeMda
ysR2QU9UsoBf/g82eeZpYgw+qJlOIzzdx5flrqJbCXp+bk2pyACQbwT5C+14rWRf
8GNTRxks87gmU6bUXVX6m/ehfBavWzG2aKO1D4tO0o0HJ0XdT4Ei4qeuL4qYfbfv
FV6m95lD5O/YkmI4GYQLfFwCamWR8d1iI6VDmwHdFJu5XsfKyB1PqQkQA/sQl+BZ
1iF0ncMJfTEC8UM2xzvdQ8B9nMEsXpDpZhQXQaunZjMRxolflbGrVK0XNnPaM/AC
goHy3EJxLN6Brn2o6HR6AnG4NoLdHdyQb/VTkAqeSKp8QJf2dYgHDBJYHw2xWhIP
clKH79TsElNKFodRjT8N2hRZNLNSRPvx49iH38zQFwd82lQ0R7EbxsaHmBAJOOz6
zrETNER1ezYH/FsuKiKzZ2RI4EvYQtNl89h6+RDFx8vXUcKE50hsIcdEiHxPbyDZ
GqtJX0rkh/CdCDqfKnpBH9lBdpsOEptaNgmZwwRiR9PLNs/MClLYKJNntmQBYRI1
D24A7JiSpXTD9cnIRsdVpuR9jFS5JvJBqXpsvTPNA8V//6pbnQQg9S4VSpHrTmAK
a+aYLFvdWNdfDuwB+EnwFUOQdF0iUCwC8nT+rtvUBUbmst02NMzE6aiwCrKcrCk5
h7kpU+1dIBWnuu6EtK4evEFsCqMaBjOoBsNz77KznzVCn2DLcNHXxCIDVn2odZuK
6PRx7w0GAL+jfEn+sgJ8vT72RdHgs68QQyfHdamWcNiDTdQorS41dq24U1y6MuRi
m7uytwTRp9ZjerIJX0qB9p4sDn/7lESrWuAuwuM5Dv+n5PnGTp/6bBa3Hww0zYi6
zmDvFhBWJGccD/hC8Owgj/bBMUXoQedq3TDgGl89o0C2/HF2CTlPO2mh/V9EtdzR
M3Ua6fQCvV877WXxUtMnPd80eFB8MDbUXMQJ3UCiyuOkknoQ1IWh5H3BpUNjJ2z6
NvLaG5kzEjVY50SYwNbJ0FDJVN5AARmKsKFTHATuc3a4E13vMhShh4z+wcXSvOtA
OqgvazW4MuAKtT+dCNU4CcaDYUpINTsJShQafQNussOFgOelqP7ZtNFuMaBcZt9m
unzsF+UGoUmNA/sBliTQlQGBipqH35Th52lLuyLKbVISUdna5Lwx2DydBv7OLGZn
kqGgqXm6cE92Ra/2DXsRWNmLMu3l1FgT6ruLo3S/x9M5L9JkpuVrg19AbUlF06u4
KIozWwLF4LYjqiPFNDtL2OONvkB7m+F/ipRE9ukStC0KqGaBAmVNYHtk8jTEwUWs
kaxKrxLnnhit4xrpq1uwVJ3vb4uIkwLl4t9h3aZkUbPHm4mbyfa6VCiGJ9jLeT5i
bKzU2udr8oPpWLgLmCjZttvRx/fDX9FbfNW+BIQjqLQdwXy7CBWJrnwLOEso/1DL
xncn1bCjbax37917tLkvAUDaN6vw3dET/tlgbKm6tq0ZA4PBN2gXQ+9l+QaJoPmA
X//SVHjfWr5s0V60YN99lafy1vkzhqQvlGn/gTW3Gas0B82OLoEgANbtCfVbXekB
G2WycIsQUkGxu53dS5ywgwNHKl7Ig8ahs31T1vv36Dgr62DGqcQA3w8bbNZJaVRB
l30JfiTyzdgYUyfpRoIZwRP30yTklgbjMlHoHYkelo7Ggq075pdCZHOocyAsnxwO
rgCaXsJoo/GZuWYWULYxSNBQ1vwHkQqh7ZO1kbXnVzPLU53xUWkBxJiRhMm0WBc1
5RC0lnWDBig8KAkAm1ukGQ==
`protect END_PROTECTED
