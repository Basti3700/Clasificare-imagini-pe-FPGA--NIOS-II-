`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nt7KPx+SwwVsxmMMgWaGbtw1cOAdzgaC8h4Efihfybsi94Is9vl/x/u/mvq8QvPA
61dvVSLB0dsdqzycibBbm0hoxyJNX3oYugYh/gXKIcYLFncLasjRMy6G88iU8P9T
F62Xo4TYKoe94QdhUY/8XoXSiAr7NkJKmvFmpiNdncPZRBUFMsPosX6tCncYtUzt
vg/5Iq7Pi1Id/F3FBrJf0OFBh+6oqpg6zQ36+uMgfqjAUyRZHG87NBDkbJPCJr51
VkzDRe+CLyi2cFkPfhVhBK874p2m9BTDCXTDFyDquhEcQCh4xQsZIpXNMve6l6Zr
AuqIt/VLpiZK1mzwgNyJtVbA2Owd7fxy8JpkUA4BaOa2L8B70c0tq7mqABHNSO9F
/myhozGQOarroeMQaKYVg7OokAwAQDcpfsQuIdrUBwn5mN4PvCUGPLOlHMDZhJ2G
LUvvio6DxuOU6VpkGM9xZXcP/H+GANL4QZPHbdMgf07M4hmWVWBUcukcv7cx/fK4
aidHDTrv07H8AyeE0iAo/MBXUduA9kGWdk+JfDD4ccHZDRFQQWQzV+U7hJ8dIH4a
7bhSgcdYR3Q+q28cSMMYRhZjVvmulO4Kj9ZgtkNZyT2qkzBVXb/XHSJBi4PCoHCe
jujD2ZP5XqtFSttDZJZvJaNamKndj6Q9kkhl17QkN293QFzXDttNXywSkTN1PgdM
PKFDXTtDPIKrt0Z6oX2cyfIX8+P+VEZwaHxkQ47MtP3LQtRDdcqnvk7Pp2/OgJc+
9RVjLBYwdxMu6eF9/xxFbm/mDFrcFRdI612GbAlAR97JyA6H5DLBv3F0H5Jbbagg
j6+865KZH/1TZ5tYffEbf7ww8ufqsl6orSIwQ/3hCBk8viSHwNR3ZEUh+cjjP0A6
BKkYpgH2THjkM0rKpp7qPIvM7FU7Ojz1k+8cTZEkQZFPF5dX/3bBx37Th+3iXMas
Ee2fhNRhtJoG4YA9RDgKWk45m1BWwTlT8xD8vukwsqNc15efx/m3YrFeS28y+bOD
s1YHk9vVmGY8ZvgdzhUhGnoxhtb/CnDMooTkaThqQQkGeqoBlN4w0KL+yaBzcn+3
lgvxWcb/vJBNsVYl1aolPuS0c+ZCHKurWLTpZ+BP4M811TTx+lSu82oEnYTbmzEc
4o46CuoRANncxwNsmJ70babJWTB/BqD3m2e3GNDaRnu5hi7Vy9mlsVw87NxtEz0N
9h0vPlPxHWXezU0W7bTCLZEjuH8gkESvkM1MXK5YrMsLuHa+tJJQkyWARkK2WzTa
4ZUvw3pca2i92ADIOVJPS4jqZWP7lJj/Ddg0JquJF75SB78I3JpYqn0GGuI9iGiH
UD1CrrKg6Yzs/x7I/ARLXw==
`protect END_PROTECTED
