`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Zv8X24MhKFp0WaEd1kYXVaOBQ3FQfCTxDGEWjtemjTpV0c+7MCXucOKmGbQx7Kp
K5e3YMeh1q4RQmo8w4xV6Pwm79+JMrUnwxWRf06kg/aXdyk/sa49HVewawNps4XB
mSgg/uKECsnJiyHMi/RJ6+HSU+U0SGgu6k0aw7eGbFqfpSoEVrk3uuRS0zNiWz2A
0rG30H6gpqIombokO7ZCla5oKcIlnXj8XPCtxyj9Tc0AlqUn0KuMpxjFYWImQtaq
YF3K1b0QEKH4MSwMLXeTYZOqAFbxhUkioXiGWnuQ7p/3W9btSWjZwzqLbwGpyhv2
p7TcGbO4KjtlYFiDVJFObncKWuD39vm253YmViB8YjbtvS+6/GjSjS0Yt5Rh975j
Mfkcwe7s1goRoKmUQGl1eBM0RjNPI2dsQkZ+7bwpD9c=
`protect END_PROTECTED
