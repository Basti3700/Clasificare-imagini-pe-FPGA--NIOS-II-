`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZvSg9+tEfB4mOhQYeLrIU5wjLkFzjzPg9620zPD2Wp3iYkm3AE7vJDw4m4WCjVNJ
7Cr2rEsGBzwaSQkWVXRsjwBkZZhxWvbvMQ8yPYCB4IA7MouNXWXm65ViHh8+XJhw
itDTHVen4bXBzcVQLYnXEJNtB1NUUkdKyj5WKzwxTlZd71gpxt9zzq0vYgGHhJJL
E+4l8O7LMphwyX16BEl2BKc3dQNWm9O4bplGh8x99pAxfTy4OLmGaDLNWVv3iSX7
LQFuqLGY+ihDWdCbvcZWTGaWbUQOU2ZmeJ2JLYQunFZH+tJd+mW0NSi/Y+3bOONO
iKNMAxWy9EqJHepArSEBzIEqSxx9s+cc6jJ8thqMJW8jpp6dEJyKFAR9mmU2SKKF
6KVPNff5zY4te5gjNW5seIOnyCrDIku5BFuWvNhDI/p1JIw8Hcybt10iWQuPXiRN
t07F6QfuH2kQnVvnVCkCP5O1QCRLa3Lyi1X/adAz6DgMMws8wQGZh7/FtWa8F75n
3/GATD94WD9VTvAYE5qSRubi88+fdaFw2tgw/ZJkxfsIq3cn5X3aR1Doqd1NGexd
XLl9SDt0w54omHUgPM20l82U5DuxF1XuQEw6WxOKsI5Um5ldyddC+ggduQGUm+HS
IUTWBYMVoEojERlU/VG+y4kEQt1pzavBJS+am2wVvDa8G56eI3nOUQFS5huSCQGH
RGEZAStjtm1KhBwk6TI4d0WiaMUnVTnvnPHsGa89Pd5M46u8xU0XTogdhtm4KRsJ
QaHvk7jhKDVc0bBaP30pT7BXGliaG+XxgffYzGAy3FNa/nHRZnzPsKMIJAGcS2nG
lawXmawKLnrY3nQtLIRDhJLBrd5FUBKImrcYXlikLZZkYjyN+UA5TWo0mRk7nUHL
+XJKyqi+2JwJSsc5H3o8QPyepTPU/oVu3qI00f9p+o49S4JZDd+fGUT2gnYURV+E
te0Npf09YP1wRel5iO7kE8mQ6zaJJKxwNKLxZ6YifTOlUuHurY8ogJkg5uGM7O4r
AXRS4+pV6Yuw6+0z0v0F1AUlZhvOZLWBv/WSYNlAZZVSGyMXd7glF8alNnxZmRzW
bPt+IPZRpoHrSSwRAc+SQogCqcBFc5iY/Z8d8krFDl8S96dF7aC2EI87w5ymbZY0
M1G3Lu97RMO2A1khR+kF/hm7HKnVB45Ll2q3WRGKX4Nf5jTHxh7Fi3IDU12GwkYd
xrFu0rIVfS/hdBM68ACgcS1KKR8s2ryuzblWvNQnj5AFCpUUypptFkIzFlWwkPx1
OuyDxyfSvzz/yiNVIG1FDRm9TE+9QZE7N8PaBu2Z04B8QwWIu8GS7NaT1AKyox9n
yNCGkJi7ziKZqv7FT2t6V36tre/97hXgHCTiNt5RjQd2O+BuUOuxbljHOQD66U+R
kHn7lbMGhNokIuo62B/UCmk2PfeHXIaYeh4fAM8NM0mc4P0X2aGBuASlL5FfYIU7
nr7VtEKcsJj3qv7EPFCORrTkx0cxlECE/PCtCM9UToetdrbwqe8foPIpYKApoZgP
s2iz0Y9FgEVX04HVSuEFK4SLwgF5fopFiHQdDRyv0Bn3xUU3Zkb0/Rbwxv042gaE
0Ky85OKUFh+DJmWR28/KcELuyVonruJyfIupkvvMM3/P3SK1ax955VQDeSiegJBk
YWcU7S5X3Izl2YBU0GfW317kMTm18pM/bpmJRGgGUEivk2eMgxHoBca4jaSO5awq
O01xAebsqbwfepgSJdsTTlsl2mJg0aygPIY05uainQB346GhrRbJbT2rtsKPIaWw
+rqYTukf8zripzDw9b/USZtylkSRidQhq/tykUNVtu5xIcvISzVVLZSuCaNE5mbD
P87Tn1sEwZlR47uUwGo6VRwIGEIGDjqifqgvo9BwwBuMUKxfZikFahVzC0aDeVwC
xXgl0MzmlLVQxEZk9xPkQSsAhGRiXaQbmTLnGHIiKr3xOE7rGXkB9WyBdePbh5nX
hiNDANCPGK3XSMfMzdjwjghdbQgtS0FhZSNwja2E8RCoR4+cRp9yemTG3WgiTKg5
PEK1jaJmzOSIkvHDUtd4ERSdUSxKHYrfQQOUmXcZ5BBB2O7/XMviwU8zVKbNTU9f
1t/H22vkoVk2Vuoo5CF+Xm2LYlxbLVXLIeze5r+lPy9iEUSitFPsFMqrEGxXpz9r
NAFJRj0p/PcG0os9yJAsMWn8h23H7I9N1dXkAJqCOzTrEONWKqkDwM4wy4USOv1W
pEvKIwxxSXEbkO7xKA4AZERuUI6FtGZIHkSCzE3FlQPMUnkDSmFOzdnV8WHTGMXp
ga+bS+h0ZnO/kwC+Cv/5SHkivmU4lusIVYgshgp+kKtYIR0KwPncG+2zgm855Ixm
M2fn4OArm78Phnki+Mq7VR9YsqXP/z2gHxaQTsKo89C2bx2rywbqMK3reHXvFaQl
gUArFG5lFEtd+oWOMCWXxxgH+6DqxaRUGvIFP16epBg7QXkO1c71ckJwUjXmXCS/
bQp5kOAVtcCpFk2PKHRxlMqZFhTTRMvsypvbUyrcuAfb0XnnwZj6GOH+iU5CxCTv
ErpxwFXRs+EFT+/e5Xg2YoU6ArcIJcN0dPF7uAgzOK2Gt/VqNypQgNCL1IZfDXjJ
lPBI4PHkk1eeCY5Hb6S14BH+ljy+f5uAgLiX31AzxhlwRgKzr/evexcY7Rouelde
REaaT2BPhfTdxZyONN4QdP6E+R1wx/nWyV6VwTjVcFGCRFWCM1gQjiG3zBdWoQtM
8iIQgkVarRW1dyXHoo+Lh+AR9Ttg5kbyz420ozRMEOtf4EbkNgMB605DfZHdaMCT
JbZMYCtLSzQshcxht9c5aMCzR1c1U0SOZSpExMuMB+T/aIVpis8YppAULKbfW1OU
VR5Qb34w883sJZuBFzoL8Vl0qMK8mhRDk56D+zF9rNuigkW14ahmKeG5Z3yQm7J4
`protect END_PROTECTED
