`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d44FWNoCHom63h74ycG7/tq+KP5aDyIO417NkdDsNeHwGUu9ri6fBrX/xW8PfxbW
E1Mu34+vB+q4ag/ehxBt/D4Cmr4CZuWP5T9djJnokZj/Rc/H+cNE/Xekj+VoHLMH
1jEjZBwdIUB+XRBUvw6168b5tHvQZtjB2KJId021q6/4ZA3siIOIDdyGt6SuBH+K
/2wmqkQtvRQ7UCrWeB6GYYbXQ3abd3i1pf2I/8gJsoiYyoe4w7CAPqxVZg92HTLg
dDYO1XYyVbrbovHxqNKIzKFMPhq+aZzNx9Io42WCrI8o/Ks3KzVl5n517jOYGmK1
9DMwq748kT3p5Yn8I5Acd7H5+Nsd+/PBciqLmUb6ylKRfVmp9T03ZcmI4AW7RHLR
DdmumFHMUcnC7pSDHapk09rDGfgUlawV+iIOQ1WbvT2IRTruGdU6opBC/TteCxwz
LKzRK7ENOR/0Y2llmOEgUTNpsRPhG/vZlgMiTK531+H29TTfL5FjbDN63fo0XHHg
yGQD3oEAzxk8VKPcv7puXVz6q41ESxcRCDzWfQb+0r5+NtzN/5q3x0TYvUGzgioI
bBGpKrhLx7eCmMsggtWsr2ZauNW4eYUjm5++vvTT0m5PuStndoS87XFNp6q69VFA
v8ZVWCcg3HdvhBjglqq+kCAQ/swK/NkuHJlzQXQEDuDl39O+aKs6KEcnPsU0DLkY
Ds9DTb5JgVu1czdODnk/suANGWjaoxITZysHpNtzWTNiqKmqi+o86XuTir/S6F6v
3PzoO7kB/v8Q1H+3UOs+nZCVAXKh3mIiSNvkYQ8CwWxyNn3JADCCmUjdyWoX1jBu
PrOY8DIapztjBL4lucm1FBT5zsEvK6KiRP7zEsP3YBPC4kC05SMfILvfRcHwNO1S
6Dh3S1K9Ykxbhs9ShP2jgD0NJHhC3pCVlO7poOkdoydJNMrJEdgqHnOwHVfMRgKY
NKr5J/bNvvG+BoE5CzUAkkVv5Kp3BfZAJCpplGLo5gus520PD/+/jThXh6H5VCR2
XTUg2wM1IHep7PkOv6vHLYhQxxyEVOgt7GDoYKAO9erDrHiR9IGmeokz33uxQom5
GdS9JEPQut8RllfFBojUAyBojHjJhMtzivqgVwooKVRLuBPBSmfJn9wvq7UNMgtN
V7n+ARs7y/Z62MACnSh7VrCFj+a1rHgJvqHExJOxpdOLAF3FmMx8cNSCd0Hef/r8
oKIVHEH+50ZisV1CzxI/PAqj197I/J3KMJ0tRylY3IBsDtL7bRXh3pRX8bavNOmQ
9WJP/VeWmqACPX29SVypen4O4sqFTmlObGOhuYPT/ieYGGSjwL+jZegdrrAdQXXt
iwxLbZKq7ofafmGlZXPenBZgHjKFXHea46Wuspu/g64VistENqYodVAapDS1qFqH
q0V7+mqISOaSGFJoTgNXfID5JuoJ3Ac47T1Lk4K2dqDLDoQV/YXeAvLFOGZAx+wX
KtNtop+nYqB2IfLEqCqz+07UNTTw3gc/B7f+7vIWi57xn8B991vomR0L0TOwl9j3
f29RKVkHeIDswxT+V1zGYua43anfYLUspmw2IKL/jmQIWod//D6wY0XIGJzA/aCL
wZnS1AGBX0+51/sVjvYBgYC0Jo/8Dd+UezY+Ah95BKzMR3jqmmoWwMPHjexIhWys
E3tDUvxCst7icMwzk4odsR03Q5T4WVeQdYgbU7Ai6mDXbDqBxu9qU3jrd6qFs+Vc
YJh0Wgvx9q2aRpvRTy6vXP2j8HJz0+yuEFhTmiVYkEXqBdYueBX1HNXW/4cmJq+r
C72Esa+uYcwbWEHD0FmUcxynHjUbQuNMAf62PLYtvyNU2mEQPf6dlcPqW03Q+0cg
bmw4QrFZkhnWqjwErxshJQHbCoFf4N/cafkXet4a6E4pSpeUlHAXzZJq+PfUkocn
+tQWq6FFe/CUnFYsR9cPTb+YD/aFKlEN7pMEPnJBDAYt41Uo/8wpTXtv1JNw3+VP
wnjeuhGBZI2jU1FP3nmLS6BOeu9tKXfZHrxNtAyqGIkrN5c1b2jXv3sJYjkvtgQM
0CoYnMxCJxIS4sP8KHYT0fvrKRtFk88DxQl/W7Lp6zBOHMgMA2B4VOAWc2yjfiq9
dRQNU1iAOZJLwGn2AHiMo37Gzx0GJrbqC4LBLeRyT1S+U4Ormelq8a5rHMpZIlkf
OHlvORJhu9w4iSirQ11a2B5rF9Wc8YP4nSdVxBuiImFuiXHV+jqRrxiDs75WtXDC
mGcFcBMy4XyOgj9KmIRIHQnEuUeHUI6Q/o7LG9cHmctvc2PGrt53fAmnvWErXiJw
YH02c71/U76T3eAiDJacaV0/PgnH7AUpmjtT6QuiHq62z4qffgIUFE9Rk68ZuS7c
PIsdCBUOhM9a8V6CoeKHjKc6hGcvO7erteZxAcWe+mAj7OADFElP194rV90+IRpQ
dMvtIpvpvt/vKvRwbkJpIeZWuT2+hC6BnhwpPsnyLJjCz46EgjrzIFcgafhpRTA2
u3LieHh7l9BXvYPqM9RRjpYxlNAWpE4+Gd61X3OaqFb96zAIkRUVwIWlBkLqnWgB
6/tZ2wFPuB7YttoULZ/SvCgbsrJ3NxJN2pUJDSfgZlqdvFl7y1pX4VYGlVwhPvFP
+pq79UY08JW5TQO65t43pKWDXEM85wZfyF664+hMNim98Nl+XDbu7fh6nPU+l8MB
CUcNPliwZ2MIo4pKxy7g2/FC0yZgMesruPO7/9ZGHNcScyL2YU7sgzWwFdc07ZxX
BU69ElFHOPAEuA30W4ucOh8OYCssMSOvSbGAd7UnEt7KvPH/6QayaYppS3ckmnV+
IwoBvgKPVVM7W28gX+PSz5qWvwp2Vz/10b9n3LtS5Q4w59iEm84J4f/yTPKS7rJ3
Dg7WWwxMQ+hfL9LtxtMRWfq7W7AMGrnXyV2y6xDQJ9iqlh9re2fmgTT0fTv8Pj8I
W+g/zYmu+ZVVh8p3lSi7+UlmyphTa2xge6w71zvvQSY1bxAL0CU+tpPWXZs1cav3
7bpzkskdjyz1hTy/wpGRlfHDE9Xe8WSfBA3dauyTz1WVxkBeOvlnSaPcH136m9YC
zO7dO6xFvAjsGu/5ZPJkaWMHW5u07k4uX9Gz9bxg+AvEKQXuZrahLsmjOObOzdH9
iK1H7mKAFNhMpXunWX8k2BpMyAmLI01MOq8lWjcsdmP7SMa0T4j8pXaFpfWnsrVj
7uWUxbsvMLTDKWJyRLtyQkpT1xDNPba8ArB3Vkda+Le1Go7tVxKGwesnRq6GsfTv
7hPzWxo8ZT5XyY31FAQ9MXU2b3Yvgd+x7UPHs6l/wDl/I0mNdiEgbdvQUwiYfvSr
+7V7tYd/W6w3bvgpzWt8zfe8rNWojYrJme5uu6fAATHNqfceDlvi/wQ1/AYc3d/E
04+4IVQ1OD64VeG7vZQM2FrNobh//h/J3yU7a5I9VFxuq7ZFd1NlHZYIQcpJnmtu
lgnIseVs8Nsz687/K8ACHDNMfUDyF1SXz8v76SnQDpKkOnv11Hsh2xkIHPIK+2D+
z6+caM1ByilnucBJz6xKbnF6WS/dZZ6WMatuU+kAJqjc0TK084z0lUFCFCfITaM4
2zzGOT4YOADo0wUqhwoAXrwN6fG+GxFaCWWTntkpvEF4JrHpan+FT+96v5vCoIS9
qQuqNxjdcoPeeopkif8U9/RXEefYsKs6pB6M9OT+xMp4mPjJnITLeHG2zyRoOcul
Olx/hf/kfl6YivMU28Qk8YlPyhtiyyHPQd3CweGbPGq10uVeXmmzyVvyRl/ddCGD
kujP+XIaW/pXhsag+ubMtVwZcchWCTJjO+F9q8VmBSrErQT9Fu91Dq+QjYEG2CQH
h1OzLD/XDt8DH6sVz60YeI1j1o8L4pfcz49sSjHvyyFmv84nuCdsQ8HlBI6qJrz4
wRxTY6c3bA26jjp6DbjxUfHrca1luj7uue5GBcTYNZXTjYLSZBCkX51mGcTKbiR9
r/hBpHkjpZ70IRUd4fETcNoXUQB2xjMDnmW7HMH3vG3qzisqXMYsDO9mH6cSQHDT
F5RIVLl5BPFOvJQuOdO0hgCYJwaktIKSVlNaehEK2m9aD+cNLjE36kZ6kS0qbKRU
AwuxQSDhEBfT8uGIZRc3t1wr6GbIHzpGeG29WqQN7OTpCupWLZcfvdpRacxZmtJN
cih3/Jn1fbIZOyX/W8iQFIsXqb/qvNPuEpBoEKwD+yQqL2cfzKO/ivznEZRwwiim
it38ulMcdl8SsAeFe9W1LrHwqIiwVcrprmP6Yt5ASxA7mMRRezBcAg0Y0Ax2wNus
U2hGUZ2sokIdZY3k0fp9sxi2oIiaeejVD0TGFHsDKgWcTJ07jpfqU0AWoRUAVpuj
S0g6Dvq0+1t9csBFhr/sH1d4AmGjzlguFmtnIWWmpzsqfvF17VMqF6+BIvjSWazX
SgJGbm6YyHilcoyF7vadcWlkr2/QaxZZeVMbFl0n88DRdgeGdWm7XL1cT9mXNLPJ
tW7K9GFtzCSJPCNNt1MBW1Zat38koIeadSvALG0SQxKDIPWhG45Z/GUySw4A258F
MeW+biz2YDufr23Cbt9Za3Zeg6oqgv9/fFDy7nq3VmZyGHc9mGZZHceVn2RoPMxE
WZsiMmu0la8+EV3dg2KD7voRdzplMz6r/V2k6tF+cVNB9lhUYsosM0rE6fLZap3p
H6W3/gcaZESA7LPTTyAuu+P/jcWOkG3dB3BslviEWcFn/EJmKUl/96uhsqRy63i6
LzNZ/6e/ew/PeT5fc/aHAXsc5ogalLlHR6q0TCMORwDa3KO9MU6xmQIGAlPue9Kc
HWqc/HAD/05kJBEzfMyfZVDv/DyFFK+sUGKtonyL98EDcXS/w3wi2Twkd3mWKgUY
GrE3skgrMqGFli+8wjovMUD4FnBdJMkr0PFJ3aWGoP/tIOdpa1XeYXlmUaRtgbwf
LOyGA9vXaIjWZpnKl12Vu/Hhxg/U2rd8EnLnePP5F/vQ/WaGXMBU9ZLomjnWpATL
Yiz5M4br4Ir7dPI1hKSxbDnlvcKb+d0IAoxbmpWmpYRPVG/TE5cSNlhs5CNJG/Vm
N1Gos0DDxfCFUK7cqt8fFg2lVs4O7bhIFmX3qM5UO3ULhCUuE3cA/1qJveZONP/h
Bn2FuI+IiRHQ9VQM5WH0Dg5u4SkQ0C1R4d7ZscQpUtMk5h7gXOMwarVo0XpIxdNt
hgXAr7LUCQ0kHzkjIPWvwZwfL14CoFTyfFd/JpOTCMwTRiLHaPXqyTbfofaet9nl
YUdIkil+MQuUFAcDrVQJaOhwnPmdEr9EMaxV8xsuUpjclbPw79d9zzQZpK1Znpzu
RlgeSJsK+T6aueSn5lhdXsvgzmAJDTXtKMSqJapc32sjfxP9Pngoptuayvlr0y/g
1QHPNH1L79mstKFkUzGkpL7wDo81b1rY8wEJhX206P2PbCgttC/Jqe6bPdQVEDOj
yy0xs1lPrIYXwCIfq2wWpySfFalcrL6OtDtl4YLjy+764ASX6BlMeXFkStZnY6vK
mdUpeYc162tm/6lxK0sFg50/c6rDj0NDWSsrRP+GrjyM3/dUTB4Wjv6zTSXATsMV
O/kRsZDN7ERUDSfA53oITC1+8gOYpHa0OoQqVD2l1xY+J8Z+7t253o19Ole94OZi
PxJKmYOVUd/5om67VFSg9LUIwLeaAEV6cIKP9P9zglXkPOyIPaL/X8hduTGPEhQc
w7rDbdqtuEbfZhbUBNbige25lVqEaV1D6VffJiceA2O5j8HXEuJZ8Hd8k3gEiELI
L2Vd5/Dm2ow/L0HbqfZKuIp5M67pt8tQ5i7syGJqFc9QiWn3ZFuag9KqDD2vylDC
4eKlZQslztRtUzW4p/2jLpJG5dB0liqe+Goo/WuaizsCKA/38ewq7Of31sYihm6Z
OiRuBsd94RTn8ZLZqSEf8H+q5onRVGerMygikpK4gzmHQN+WpJrLzTsahexJyGs9
eH2sxXrvxKg3USAr1rcUDR78V6MYBI6bV6QCtViL2P7Gb2+MzMh1mImhF9xDq/Wy
X5TqbbZsSftNresGvpxQvmI6PAtnnEM/W2rW9y7UQarcguluAlKzgSePlM0wbl1G
Hp9D6QPWFMI8Hvfuu3xrkHj2UqjPU6j7ogu8kqueuP5Y9LSC/yRi7o97ArqYcgLG
r9OfYswnTgeREFL08PuOLYS2VzJSOQYeO2eXe1BU0YcNCyEeyHOFugLmTeaVZlz9
GKgDbpfdQNKv9K8s5sXneqzbod7kfBk0PtS47s9oXbOXn6Hat8G7YctMQ1l9Yn3d
OM4QpfuGq8U+AtBk5Muhrk3j1Crps2yBSO3Rmulbt5hl3Yhoq9/MHhWhMaXzmr1X
YZbNgj2nt8x22S3h+wmzdOM9dvR8nPp1VmT2l2aheSVClJ0LR/yyLkOxR6ta4JcW
rJ1aBG3YP8GeJLo3xyASv4ZXBmffLVvSCbYEoRKXadj1L+DdMYNyUR8TPGGBVSNy
GVPD9s+c4JswsBqgeK3MohyD90y6PSv1zATtC1xI6UgqLH+P7S8+UyqN1KsxM8Gw
avwWPReNVFd5GslsWGCsWL8KOM0/1QLJm1vTCQx3REgd5+C2f1PU9nUnXlxtqTFH
jxNGgy4fb4hmAcjCNt+aRCDG4X8s2eqzGCMtcIuZzzLFpzR4j+3lB1aJr3ZGEqZe
wEWcffYU3nxeBkHl8V6iOImX1+GM95GvSh/AgGzOIVVx3e4IlDqK7/jD+S2k2vjJ
yUwczdwhNedQhex77hrXZjlNYG5MdmCmRaTOg2M5Ab4=
`protect END_PROTECTED
