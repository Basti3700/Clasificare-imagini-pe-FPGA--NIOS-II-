`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8ZpKA6Mbt6kcW06BBORnqxZ6bZgjdZYgHdF1URE7eAwlTjHP3iSzy9J3sXfujCy
1p6SaWvmdT6wZDOi1qDyR2QKBxYNq+W2ZIqYo/iUkbOkO0ULTkR70H1GVXfTQ/sy
IeAFwEy6TSDpmgErmggJ/6EbAn1lHw8es0AL9xownwKts6d3QKWyz8KqO2VLKyjI
bX7yTTeU8xhlzGLywERdWeqNjPsfYz17/J691P2T0s4b1SV0BGb152u9Md1bMoEr
Feyj6DInr4S7S9WBFC5piQMmwVX83zS8qn3qfzOHy3uFaw6+U/+GvZ+ES2+5fd8G
jw96uftRAXOicw5FQ7B7B6OId7ZBgJETuLxRZEkc0HC/uEvbw1PsC6tPhp2Wd3ml
xMOMBjw3m/eWVyKAUyfGps6xDIio7VuTEy/iu3EplQlUJD5cmYWLw9gqyv8YlU2H
4un4F5nIPFWQOCpXyhDYL4jypWnOrcTLE0xi3PO9LqKxU4OWM48rAMWdhfMDNeeS
r73OKSak/H4iugH6AxxqIVhXY+70667n41fsCv45hm/n4t6bb7m6WwNzDNepcjiC
+S2jOwZTE8HLlzwyvPGQqG/rXX4wTYzAi+AKEVgEqnVYkRUdraX+fYlNjLe8fGVD
I56WIWCJXff68KeHXwm+gvxl55JjdQHm2cs1QpWTS9gK3tqkRKsZMMpkmIrrsmLs
eKN9SxAAIdgn1kpQ4mqR8cLZMNcKVegV2PBCl0jQoelPpxhmHrpAC+ZxsJosSLMu
cSH9j+IJeuKH47Ofv1H8zG3Th274sMbapcfoyve+fmz3RqFM3g8nutTkLiENhvWu
LibBN8e/DLome1/sYbsDiB/e4uKqrsMWQiaDuonWbj+rHPVMYxddxfkUHRnnx7as
V+oSfuN/Er11HEBQeoGCl0TbdxeqDcUjuW8GeKOXKvVlG8sDUg30KYXq3XPvs3Ra
njo8/AHtxpb+mcGOYxirKNsOB71/dQIdIBbojYrDPvUwOwa9srnbipRIPGkMMiAV
8yFfOO1CnKWWWVkQuqiXHxU3TtiC0vrSP23f6wXZ0M9rslXnu1wyjvMzDBrxafhU
Ze2OmxNDfWCdIlJbUPxd1dm19uTXsw0BsWFFFBdWkklnVRJb6dnaJ2p0iWwC++2g
jqVbkP/EjvhajjZEf/I3YxjbojnY+bFQjJd9SUJCUl8vHI+2CmWUDBYspqWEmj+r
oFj2gLT1ftTFP2HiaflbIeVZtC+hh0v4ch5JznwAOriei3ff3IS0HcFTRfvA6Bfj
2XeMlCprWMaTzcXB7X4r2AqkRdIHkV/1XrUq6m6M3I75kHx3Ak+v0I5QXGYRS8gK
OH0Px5LL6OSbhZbxxFWMrtpHjAfcR//CVjBf1vKK7eBrzArxnE3/MdKoIWA6CwPK
e5D4aVXmQ0h9wpo8Il/1FRQ+GhcN3FSngJWVoiw1oe5sdispkvvZe13Gd62REsCF
70dUxbA8+GI9USK76u5RE9G5lIkpDfJV+IH44RqeQnX8fLVtARGp12MXkC82XNQG
RQRuDbx4gkUSiCgW6DJHoV3M/gRyankdLmYKkax9+4Qz/LWyEVGxCIPcsybSh+qb
FoxRKlOpZbnmjNzBgrcpGlhD6s1pw2B2jT9kgZFsue5eBTBzowtfdYKJg/Cz1lnk
ufF2bPwtXaYrbq1LhroWncep81AhQi8QvIEnv1hRTTblSQFJnbU/wrH8G0YlCUyN
jAet1KHKecS9VX0/+c64Yjr3efGJy14RnYCbiIl01PR2FmGGkgUmUa7mGmVfMTWb
tXZK8BvpdblD1lGBMVoGrvFyDHX9MxLlYK+M8JuknMveLE1F7Nlg5DmbmlN2Q1oe
c0wAwXZu9O1581QN/jjuUmZLsmF3g8D573t7B47OU9nvLRmMivKNwBqRjAPiOUX2
2JfTmW60Ca/o5SeFEojDCSx1LTAuAOgRF7E0I2OpWcm5ioKVSULBJOui31z9DIAp
0k3d7MYmOwS0WZ8a10ASocPd2cJLmt2AQFp4rF8GpOcOQzwQQ4tf8fhk3RWk8Fn6
HU4oVCGWHiAJezdY+Ch4dGtL+lcMcVv8IxXA2O45uRQ=
`protect END_PROTECTED
