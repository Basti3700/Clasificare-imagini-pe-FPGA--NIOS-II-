`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5zEuSdqj+Yqeuj/op6edDFdyvBPyNQSzmJxMyHNCnsIew1Pa61NytPrscqcamVW
GyIy2LwqsOrkVCOGcHfiWwT6wZbW6EgzR3vw7VnCgpPxG64jG51rQqtsYfqNJrsP
YziJ5FFvL/Nx3zBa9njZPrclG/P6DpzX5JnN6f7S7pFUnsqIR3ntFr2MHqQghG/1
Ahl/VlyyHdx77eheZigmADFe0zgdvcI6Uq8EKpXpJ34UdceGYUBzkuhktWPROYNP
kj9pcr2gu0cbuvOQfm2uNhCmg4dz9ZvTmhaSVTlGu3O3/DOdjvSS2H9PhoPvpnT6
ayWi6NrQ744emv1nbH1xUY/46+klgVvGvI6PyUV9h1H00/JiZerlvDfq27E+NfET
51eDLrQFmcq1c8hWB9Rya7+5rBLYomnvYEuai1i2Op+TGFDxvx9f3NnIvSAcPv92
s0+CRTzLogVL0QBvEq9he7Cp3QNyXWYWNdLKqDok0ZkOHe155UCb4pZVuTXsDoHX
`protect END_PROTECTED
