`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkxufujoNZ1kdkUZaqF3lOtWoYcv0HlVwaaRfjFrcLUSRdsJgUiUhA/xz0yBCmHJ
M1KE8rQiOtZ3a7sUnvJ4QoDynThqT0db9ESC+X2KQGLFGeg8fVlTgV55wEfyw3n0
DLjb1BukIXPyd0274mCjN5lLVxDwkHlYGu48vzTeb9ckWI4hV0DrskdJ5iXb/AF0
Jx8X9/c48zAZ6cRz3MHHGMT4fx8frEwaAovYaYO6C+gz+Bj9pLPzd2EFYbaYmbRp
aQN5Mqy2j+Ey7X607jkt+3zoHyfH8dRYdZZgxOHg8ExuyqDsleyzIV7ZpPvunIge
uMkVve3nPU9blkKwWSO8gsqO9Y3x3E+zcDFizTL8xtMoEXEutd31K6MZ7G8WuxHT
`protect END_PROTECTED
