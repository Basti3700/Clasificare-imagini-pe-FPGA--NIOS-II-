`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4gJR0LHO5+EEIEjZy9h1XT3UM+X6FkmWZdhWH5I1upJXwXwH/s8cu4dJ3ioSOa0
lWLIdVua6kiJxX8EEW1D4IRx1kgMvvbV+RWTI7GzfjOAF18kX3UlzBzToUqmylvK
UV7Zax4chB2VNo245az6V2BUbbzJkJRn6C4tWJTjn73sdtffsLR/retaqutP27gh
P6Vs93I84MJLcBl9fJYu0th16VurbRJWtRLJTgnHcslscudlRYFJkLuD+rsf8LRB
n1T5zL3k2Ka2ghN4YAZopf6+jDKkfPl0C+oaVrWBC31bGzFiZmVlfd5KcM1LVO1Y
pxi+PhSRTm986gp7cKiM/wvMt6FrhIAtIg0JMFzzCmPcCH2x/BxNlTX+L7V6q56u
wNv1TSi4OVy9hhG5aMy2bt7ALiarTiBhC+fSNd7LiLLgp3bmYkNvJhppxDo0OyVm
MWloivNTOmgJJshtIRfyR8+3eBitS8wHymuMLuucvQ3jTbctZa187O+S8OBPzV6h
K//bv3K3r3llMxRiANBqrshCD7/Ad11flKzRcsWARA+1QqQoWM0GRwW+p4fd+qDo
nrZkVNrZRgoBnqFh9OnS0A==
`protect END_PROTECTED
