`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8yg77QfK3H6q9fC8JWHhtZjx2tbx6ZsT9SMeQODYQa1v25iBBsav5c7GFCwLHI0X
3LJyC3XhEQH4X5XaWUXfpcuvhSgYPCGGOuG2CcMTKwV186U8ZroO0GFWm4WJ/LUb
0CxlwOz5pSuYcQT/dybXRC/AE/gHx46Xe8pGghGnRZhc14IqDToCPQ2zROleS0fK
tXjGKFsYSaEvUY88/1/SkxvcwpgXSy5g6EY1JwO/U29+uUgs8mjp2p/vXZ5KJiom
zSY8Tq0hXEX05in7Fp9GcbYLD4njWeBwbkzIrhgol064Hr8pxwqff2Y7yn3GPh4H
9iAewZRACo6T85G5rQr9WdeKMy1uD3OWCs52pIbqDHbtTXw3t7KhmEI/MQkWe6CL
29fDgldDZo1GsvEfMgcYd9ZAJ+No+Itk3S5utNbe9xyzI1FQoltvnnq2OsivHVWV
kn3+nKa2utCnMfcCZ4WHncO4W+XtONQa5i3bmjm9yH6LqifATSIVFa8Bl7maxamd
BB5j3h50D7ib0PgpUAVAAFK9DXvHxPjbr++1queC7xAkJum6xcI2uNx0n6RnkhAQ
09rQgyCK2/fdvwePgJWw0wt+JdPuDwKgXCLTQ7p+tWF31+47PKeyjHRxkkHDDB0B
kHcvRX/WKWC2nQvHKp7Iy1xpEc1245n4l6O09XP34064theUaqMJgJUV14afn3pn
LXUoYPmoX0p1LuKwvIJt+ouPZCp289i4IKRH/zpMiUemry/OJpNHnpxvRoFCa33w
/RPL/dge/afHIRjfazc6sPHrk3FqiBs39elmD3zxTj1qFAhbtNW0z2on68mSd/le
af+LvhJEtAk6rRWfNi5RsXfr8iVv9BpYJ/akAeATwbR2+a49ZmFPdXleyOQ6jWYS
h++MgBET1zUxM54YlgBOdLtOn+jEU4Bj1u9aY3AnMEwVPxR2IubaHZC8Fwc9MHNI
oy9+0XG35D+PHE3Fmg08KRhOhWg4fSQWQq1TdxjJx/2rFkV/f/sVK2RusPic+VsH
+nRaoXo0s/c/poCgKf/XK/qU+hbclO0BSZg+o5a9dVUgg4KvVIqsGPH7KKGg1KKA
tdP+0pQ6Lo0baY2XDn52r6PNL8dgLnBBXTMTLeHe5YEWnJYRjggM+Z8rIJV5QaI1
fUo0wmmFr98dzTYiNX2Kn5rw99lAMPnb/UXCPhQxKhIPjaNFXhuPhiihGwPfe+wR
cVpoZZhVUsi6ASQ6q00fEtXaNuJGKQrOIdqQPv4/LLaJCxXcjLYsRPoFe06ctg1U
5IBarRojWNwlarc6V9lMxM6bgPO/7f6IW0nw/GxGaCjLuL8TXQGf0f/PtzCukyk5
xr6Jjavl7dbPL64kyHCv0sAI4n9YJxt8KtGMurRLdG8Ebag9cOGNiDDrTYn1jpAV
iJP6g00vYGfcZatyJVDKgGHSPK9cUUFmT4rvBGVyBwiHU/kfHWzrSRg0y43m/q+U
jI7URxrUB3iZZ59KNTnmLowv3mrpWJDiFUMe6BBeoHQQURs2UdRq674V7HMdWG7m
KhvEBafZ4stI7JFEyxQMPMz0R+ExUEfUzkfKqyi3xiWMJYHlwIwL4Ggba60POU7/
Vx/2NHtOeFFrzT/AonDOjQP1LeQ1/2iHi3dCA2eYslS+JLn/mOojiDaWOr5ehIWw
97ce8XGi3lJql17vcvAbmF3+rAL0a1WY+uu+6uO6S5vLO8DYwnqY0Ao3hedAwyth
txl51wXUe+BKPQrpnvICjQiPS3v5rxA0KtUido7N6i02MQ7IP0j6MDPxODG6Ke3U
GQawqF6DSpZcNnD+N7bjY99yDFpxOX6rQ+kL9zwKqLnoojA3OI5OtQkMn0jWqALA
6teG8uGMo3ee9bXt/uprOwAwQuC/v4W5fxyFHC/9nnDMm1F9cZnsy/kus0m0mMTr
vBclJqD9//6vqJc8upMCQ5wF8dI07kiKeLTlFlqyy32VGvKyMXkjJs3/RudNWybF
wQ2Bkg+zMxUMcRydsROUNZKY5lrTSz8WGnLbt8nvevQ4+bVJOJ7JXxqo7xAjcv8I
Cd2r0ltZaalsDQPicFSKcZYJckOa6ojyWNlepcapKPBXMPDYBQ4PmMLXjOChRQAR
1hs4c1Usd0/1p5plFX/uTzDPhEgDLUF8W85iLy8SNPoXPHn4WeqIE0nFGVT/6swT
NfQBOqG3QpHGWjGe29BdPlZeyeC5rjKVUn4rSxnvPu5HnWftRAGBqTayGEm8VC6F
Gu9Kh1mwxe8xFhySFBceIQsDP3oB6+kwSdG0d54fzQ4RuNh3eVWUcDiKxO/FOjXF
glIdIKIylWupQry7a3F/PxkXPQD8QW58yX9NKfs8WzMdwo5HNu6BL26RLFQ52gej
fTlWYJFC3pPybUkDYudk0+yVlwVrXvHvVaJrX0y7K6W+zVh85DQW4VEE4gm25ujP
3oUCMLQADrbZiW7IUnLncHbfCroW1dGXGjBudKpZG59LnCRiSsUHCjCQUGVNdhDT
v8zPf3YKanVqpXNKB65fuiRSWrwBN16WMaMLE/38LSKH56oPdKzNDbii4z5vHM9c
3L5ELetKfbCZ14srhY2/ZyQRcYmqeHkF9Mf8Ui3ADD61mZpNo+mk6YQQ8YcIMLqM
twNjgA1iAWG47ebT1ZPNTjEQxsBVoLC5n0AXYGspPqBSb/EohU48fCh3duHnK8xp
vOuyMMJrgX7Gz2xWERTdsfjTNw3o7CcRHMjjnquCHnry4lwgg/Iuw/oS2e/dfbXA
2WkQbPkV4q94lxFQMdW4Jih0ZwRWE7g5sPslRf5Mg3KtWuap9q00NDVCTVxGw+iQ
iBzUMQ//68ONX4j4tYAu7XcYKgiaZUa/uNB9JZuoohJExR088HwWzt5Ye0bxtxrl
5aRmGn+GMyONYySZbgn81tW8Q3oqaH5/GOFI4paiHPvLX0JkO7hHT88j9pqHwzAj
bUzsWSLID758nkV2IxPl9FwI68gpdFc3sLCbCdNVWQUwcU2GGrFgSMVJXldZoVeM
yffdntHcaZ50B22llJMR7muvBiJV86jBWpAZ11LNN7odTgesgDzL2HbjqQmmCf6m
MbC2GDDfVttCYLoPr8lxyH0Gy9GZjJH6rVKP8tvXLpDQ4YhAOyWRng29KfZqqSBc
5EkgchtjjPegNym+eVNRX4eGyZAXHrhMjIF7IsommbBiEUucyMbciwuciiyYn1Yn
A5JYaW1YKzDpGDT8kZlbCzNLbf8dzCzTIYJ94baLykL5YgPlJ2ZUToynr3XvN6yx
bJ+EaqxSf7grSwPmCwl7sE1FYWichEgbwqYjGROK2dde7wu78OxKFwwdJbhxcfRq
67GccbVczFCTktcWw9/N2RwZHM7Q0mxtBqQ79fbx89oYPvga/uELXeG7trfXBWFq
f8HxT6yNoPj3VoS+2m22dFOGBD97EVGkBFKQ/1YRt0Td+C0rcjsq1QvOS2OUC1N0
pP6axYO0UoghmV5Su6VkeX/TVB/v7rXhBxH/Vs/QSrLFXWzCSHbKXyYXIFnMlCmL
kAS9oGY/DqXyH0wkRPSzq7dG6StPdtx4rO38IPl5kbJSe0qoG0RYv2KT4uCjiDPJ
iojLr1adwWNR/fz6jpdWcKqmtdnUAQATYEyMkAxMS+8MQBIgLcfUQA+Kz6U00W8z
aw3B1MuhzC1L/1xtk5AIT+6NQ5V+GnSKdzUA+yroU2gVC0m1IslL69syixYqL5lG
wgew+CwzhBwzPe+px18HhvfE9Tot0ijCzInsHNF071HrDicckxqlfCI6WgbtqmSa
B0UMX2z/w+5lYWO9y9VnBDnXr8BlFWWjE28NiWzcXmQtRBXi8HBVRkzOU++/RfvH
WYu7A1TfUUok38qGXNbZOprXQ1+KasCtNkHFcq2fBVT/ZlNzFuA+59ybUg8WTE/7
nhuSnDB7lgigWXX8WlgOHAJ2Yd2VhT6xJ0ATenHZSyszpfjD4dIZ8jxUtYJvt4IA
Am+HVSl1jbz5yRky7D5+Wf1thyLIIEH6b9gynQ4wIsYTJU3spE2TZgdWX7cp0E3Q
Zn893/d51rGieYgCshpAgYMBX587ryFTb4d+OXDhBMfge97d+Po1JD8w8TUZFKVP
UaXHpeW0zYwOeG18BQbWHU+0WpJKylLJxwrEUChIQ17A2L12XlQC6aKtMdtFFQEq
QpbOSL13VJ6jWrTK/2gfbtPdswmqzb87/lfNAbrDOEI0X0zM3GMkd8r/dXiSsSXs
mYD5XOkCuTpiCp2Rxna2pDr3dlBeWMmNmafdUh+J2kYnNToHftq/vIfesQzIxWLJ
OPpWZUcpLoOrnVNrSNpq+xD6JhRekSPHyGBp81hdpYxvTFHMKwf+hdy9XnqgGcAy
yGvH2sUolBvM14KJGKn4FS0HmOV0/8tyxBGon46Mn0aI1YLXX10Rsmn9Wbnah7bq
DOsXwlMx491oeX66u9wmtfIZHfRMLMHsFHXk726Z0PvAa9EpytdI1X3vH3SCwTLA
ZkF2ED0nMq9PIRXqTHGTAvIesr/6rSDwTQmtVfG6yjSzIBH9GMNJQ5jFd7DNGvrr
qLeB5zwLv0bTBwUlbFrxcLz6brssR2oxU8pcdbqbtXCFDTJxCj/z8CXIrexp7IMp
8LjA/8a5HKollv6GD1/rlmSmc0QR5ePTmd/gvSeiYFzRR9E8Cr8YwoRoA/nFrzgB
o+F2J3G052jvzBGGQ5dt9WGMBqQq97v0xAZfMnkqs6xd2ttNVaQCQ5PLMgpm/+ZF
dZBuygcd8bzVhKgBjoWugutKqIF1lGANi7FE8IpkNkWPMojFb9KbIbsSeokDuN1K
swcDdOzu34/vyHIe7Iyu+qXKosHszuG5MEyNUcXNJ1oAwE4UnF+F3zfoaI87kNo6
feOt0hsWc1FEuWWMRLuTfO58SjDKB+9bad00PNa6MSMmgripDgWs6dcZOgwY3Kpi
xJgg8nD8+H6UY+2NZ4nArvGt5rL911E9z53/3uORFTye6+ZsNnfK+3h7jvH2aJYv
8U1abE8S6+W2LDic5DWu3T7EyGlYYT/NrSZpphM4RoUIj0DsHClxM/lhrO2vrwhh
ncEwQu4+4/kfhdzqBH8bc3tgpXSft1NQ8gYv2P6IQS9CP482+jCKbgaJpVa0E6KK
LcHg+NdEunV528KJeoJ6P48ohcd+PBrEh7U42RJwYvh5+TP/n+2PEUsdOJzthzBt
aJPvLWAsjhFf75zhlWERXHnBlGs4Sx0tVMcxdjcU/hKnboG0Da8SrPPlks90g8A2
DrBejlBcPp7CKZMpeqPdfxybdyOmo0UCIgggbyuWFu3lmD7MfTir2vMFI5NEAmO1
I5TMy7e5pNPsqacp4vVKFwY4+eY2esLM3xLsXHGggDk921lNw4VNSzppKxVuO9jk
gFfRJq6jev5HsDvint/yw6DolKug+6TDTEHIUb/Yt5tNR9lvwIZpR6xUPaBdJIFV
ITj+el00GAEw3CLmRL7xPCNF2tHH4qHf2ghejHd/78WGw54ihpO97sUjc2apP0hG
9HqOxu+d4amj8dJy1eMiDyvJavwDKjHxQFJZzNgnBZmpWNwD7Ji5ii6CjX1WqTkl
3HMkjt2ECJzm3r1fEiUdmGWpmnF6v7nL7Fw+HUvtsAwh2ixu5GWtRnPRddujjvaF
uf3WayiCeFceXliP3WUWbIqzjthdoldJGl4TXMOmUIzsLoWD2B/uBxPJl/MpIvBN
i6wHdCAgElQ1yswN+hWiUXbaCkqcow2nTzWZqKF2axJp4ub7I/HXhOF9Qi4ZWj8x
J1w10TNC6QLauMOz9yP/QM4nCfoYcRbUWj7Rym2Y2D5K7VuElyR8qKWegUBM4IF/
BaLNeUMnu33tIMtDsgdGTalI00MwpRGZ/68yhDMxz6oARQXjGnMw7mJVoSQC/3Y/
pjuJdzuAFWa5nJFBGVb35vqk7T3Rg5LVJt5U6Y0c7eXNLqNPDGA2lEG0YUQjposN
db9HsFDnFxwtA1n0c/zOxLXZm4n+jkMZE7F1g7FB6P2k4dbtxHtWIHXnc2YCaR/8
oD7AS/LHIAf4yaWlkICYry5ak0jzY87bpzHrvWQs1/GhoFULeFmWBYfYChkaQy/t
LhknWkGEfOsbpEb/S74zIeChKWz6JjPvhre2s+QtuiZrjhSQBB2X7h32qP3+q+M8
tGfqK9VQcCskklOLTSg8+nYbPd22MAEz/YkWxUc5mBhfdkVGOypLow+YPFIIJCC9
NlsmEVAKujGHKM+6jh6ZjZFBLS/ZD8aYtLwR+XjU66SJ5c5o/SE8J2Wo0cKUZSTu
+32Xk7f4kRsvzXP2gyCbnOGeLXVvc0THW1Gk8dxGL/4jeOJKoYla270yeZjSyXJ3
cwsv5ksCvMtJHjdRcll6qpLBfE59KhYvbZYgTN34TqccvXliRxEHGjSYeuf51jFh
IHJrC0EEgKyrchQkQjnLgXEIy3Mr4n7GNYVvsOBsrQTQKyE1sgr29/2DgqsS7Kgb
VTqVr6pUzxO1YcAb56pper6rwyOzi1zeSvQIuNrZe/t6VII8NhuKo7/Z2UK+kX31
L2TT6cj8WReykjXhHnYmnNpyS0C59ooyVEOFLPNgiADnGf98cPqrCb/rMsbgq+3C
HDO9eBDZ7s96pEB+JsBN4F0aUOuvQASnEgc0ZmflcPoWydx40PkAwPWenqwXIeWo
GdgyUdiTz3hL8+5d+ULOXSzze/EXQlMdYzL8d+to89OcRLPg8luUvMbl4AVa6nGd
TtozQ6emxRsFP1XmE/uWuOEStHT/wo+AsDYS6YHVs8sZoNB9SLZD08EwuTBY++Vq
C2qOucuzQLHUwkUsAZGEiGjpmRWkgxgZbcAQZGIFOxW2iftLVzUIMk9QnJ5LGM1R
By3SC5kIVEzEZDHdl+4koWURrNpODdPXWHe0x7Qnc/YbrAamleC6RWKQkfSSFkEA
lUi0bxar/qrwiWeSTQUqpyWmrGN70wb9yfwf6EVH0EJTJY0sWx+N3JiVzc3DgaMc
Q2Rmy7/mUa5wsuekepeKbjJYJvFXrX/0USu+6MZ55NJfZGrUvaaM6OpK9DQSWlpx
hU+GWdx2W/sn7ClWI/E8FE0RfKOw/A+hestROUWov77GQXq4DZp0WT5EJutusXDn
Rx+vXd2ziKOzY6+qbDV+hzLYf/BgkYCHhrxcdPWg49dg+tZaPGGxuCTg1rrDMEeO
+d9rl3Y8//R8nturXqlINobd+cPBlyOav6NikYIxdCysAbc4BOSBOysQKZtfPxy3
FrpMzaqjnpPM0k++o4Qtb5d1EKLyRgoLJyv2bj1s1aQ0Nw/63OLJHKlUFTOtdcFk
ZFtRtbDPzwr8QvgFCMTjB+d/nH4X55itxgxSMoYd0rHGjWyMyzmYO5BzMPgblkfK
0nAylzaRrOsb1dhR3cQDH+SR+bSvTgxMsqnNTc+MLUDqPqhPPwL/DK0v9GCg8ysK
3fpz7wU7maem6rPjC0nTaxttlE8Rhz4cb71oOaIbkgloE0/hfo3dz//AHNTidTOS
i8yXPE8y+IxPuTqnCVH6Tm4fi99kSEAENDlsAae42+G2z7TXtBD8Wgs/dmoSCiAu
s7gQsY/ubVfFNCEhegSq+ixtSSsAXsWw2QOF1aU13rzLcIUUBtty0Wja+vgoc5WV
+7CyIy+aBmDJP72LFeiaLiQ3tI/wFJvMUvkFHSkDbP+ecXAUCZQU6IoLoGTaTRPx
2UXoSpxUxWJaLNDFrPaGRzxBYvVnZqqBYgDiAKKdS70LRabd9fmlIUpJBq6ofUYo
NWtPtFu3oxUIlz56ARBJGRei0cS3fitZIVUX6zVkXSPQWQqAtjW+nNPcVEtfbQLe
Gjbeswewnihq1pA3WLGmJlezsgE/t5DAUWE1/s8TbfkQyEV8eBvWTAIcYou7Qp5/
g48ZEljlCVFjFP6H8PT4Wvz+1wij9NnI9exycmPRIf0nytTu3KqIdJX7Wb396TMg
OUUxHbpNtBsmKIiyucMB6KuKMBXkNfpQ63PesrOIf4iuNeLhEIWKRGpBpV/ebK1m
xFT+HP0R0nWxHwzaDfK+AHBhJJ4mRAhU4/UcCYH+du4x+mxvYK7JJX7mQa9SoN/k
LAmZON4p/oRLFvlJ3ZRJ1GjFKDg+asBeL0vbSwC6pIF38F1pjZFAvEKW+hQ1NBWY
1YdtDdROtPGEz0lvWPOS2KXYM+ZKiQrhhclbEflnqikmfmIwByXcmgKrdUYVw8cO
3ZJ8B2fWoLD3cTDOqg/jHAsKxmC4oFEHreRR/+UwnQ1BZmk026Pyro3VAq8vpVBZ
dUbtcpYR9inqD2GojY1c/y87UH8k1GkhC4VzlynZl+NsgpCpHLF9lSQUl/McYUCX
xYaVvl4PozieRsdiuErtuhchBb5RvJZwbCatO/V7u3MYmQJgp8wDSqaBEo28fXzh
ezFZD2qetYjABR8tXupXMijQ5CM6klkvf8jUlEP3N2a6ZDg6U3diEtmxZXbxcwlr
UdQKnuNCAdUGxmelXLXIHGq2kMQYDIe6Rt4H685UZpWG8qqu76Rr1eCnrs3K/dzk
Zg1z30vz1ZiLS5ZjGuGOsCNWCOmWJVc7SJBq/urEBQzT4+bcqsJ2ihAR+1BA2if1
/awG/ChYFSGZpTuxBk+J39rE4SnHdNEBcYTz3Vv3U75VGfh3nMuoBBdoxCbr5+k8
WpqgkQwrC6Rf5ZMCYvMenlDpuFPi1f/0TdaMJDpRAzoVzXPaLHUYSq66taoF3tV3
2zjwrNOMJtGfLsJGXmaNMIzBUxtgCa85EhQOE4Kj1JZAsFV6XBR+2Bl69jjisRiw
M4CjM6Z3t9DPDtxpB6GPtlKB0+fqddjvHLNcrGRyMMg0JeihEHYpzbmzDXEKQ22G
uhjzgWq5wDPZF+On+hQK7LiiK/sx5gl4E5SnZyk2xyETotMz6UDzm02VwKLk5s7d
GLc8V3wU1WY07qM3K+DlwFRC1hkktiziy9BE0c/Njq8lmWAl5FSkfKELBX25r/Q9
QiACMbgM8z3Wt08FLp2a7G4fQ7ko1l1FWNIBvnluxZg3HBZk2NtLKK/ZpFv83KPY
QY53R4UR3EpbQSEXgD1iTw==
`protect END_PROTECTED
