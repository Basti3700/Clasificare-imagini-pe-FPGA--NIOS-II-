library verilog;
use verilog.vl_types.all;
entity fiftyfivenm_controller is
    port(
        nconfigcore     : in     vl_logic
    );
end fiftyfivenm_controller;
