`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zdIyVbpO/QMrUFLyTD/KkGo8iRUAcvB0IVux+lqtsuEdFmakpWK/Nz5xNlKeS1R
anjDTkM9t+aAvJ9rgM4BDoYb14YLWkHQvI4I0E3xhpS7NlVTf/to5HsyNsHhhNSl
oGIX6QZw4JsaSEkGpfwqBvdoZmAVC5Rahm+8iyewNY1tlBWj8PPKsb7gJc3XwBqD
88HvjhnoXZ3D++dWH3SEBzGb5IqBUTeOI9Ywg1jbDegSEDCnMwPar2ZJgeStTl+i
dLCw98p86LuKfeUFGLWgSqkp8CSDQXuE9IaWEZmNbD2APginPdHgwDgwvlYvWTNS
5+ENVeziXVsl8ICjEolZZLxxjdznozoY/7Wc+JBnpfaFS8S3ZGEbmvg1Lzz0QlDP
zuYL0xNedZmKmBkQpadETpQCl0NZXZpqJOgslfLOmS8CgYuIOoNRIEV7nfmtw+mD
SWG4mczDbhCIeg4KYK+aG7rlqD4Qzv/sFIcMW5IsVF7oEZ2NstslEmp3x7g0VuUu
`protect END_PROTECTED
