`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cMMcqmxNAyCgT29jEZ/zVcM0cqQLaf111CXIo7T7QPk+zONMzvj4QJLGOt1nsNST
ATvxWmhbY1wZBnYRA0YvO+moMD81UsjTl4drsLyMfOZNPMfCbMmrPgzmgvU876Y4
ed/xrfipUjMlXS9Wotd64A8NvaKuB/aEHIWY//qRSZbGwux19ncpFOjKOtKqbNIM
+aq4PwTeg6lcK+YIaaYzoZ1w3pYYBf5kr+JdvDRZbjCdJiRh9ymFS7xc9jmjyUX7
TmRX+fMxed5Xgxuwvu2YCLkUUz79V0VHF9QNknqbyxI1okeUw7CfPOcRKic4EGqE
kJU4sD3pF5QbhyQHd3unjFfZzQf4SqTP/cL8QFjA3+wxXx2gdMmjEjKEXE82mfkT
YkL9Ys0dQsvNJWDfsVcsMJoM5WZkvPU9DluS2dSsxjC04j3Wa4y3DtfQ+5q7tEJ7
eCGkCfAKi7SIjy8ujjGxn4mJsM7iEyLG4uWW2/NysNOaHwqpJY/mNQPy0yNlhA0V
791A1h1MjZIscw9knn32bz2y+Z6DQaWM4NPQaQ/Jyu75K31Owpro22ydoZ9JJxbR
jq0iMcVEu/31LRRlPuOMuQ1ac2tt9858tQGZ8n+Ldb6hIBQv3hQ7PfbcEJpR4w54
`protect END_PROTECTED
