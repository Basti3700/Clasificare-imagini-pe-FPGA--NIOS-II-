`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrHGZMatXyv+Ra1OEpRCnthdS/IAjaFNHPS4RuKazNtaaDLPBMD71hgyPVJgnTgs
DIxnRcysn12PLKE6w+C7TazsdVmRUJ0b9lam9HL57nveRDJS87HzidTIUk69pcuj
L/5OPIyTuXKdY7Xs363EDdytUYas+ObzRkwpOcHuliKzWyjBWJJefwuzmNowiKNX
pTgwdUY8AiCfzSNJM35iOljMykAFf7OkSQvYtZcfpWxDe+SvyeI6N6pjhv2l6eup
/OkCADQN6mELxq81wab337W/oipDvyfGXItZ/A2O+nFY7MP+o2OvGPw6CSaS2zOY
CYr6ByTN9HtqaF5Oby7zeNeTIYF31ohWbP0RNCBYher1QYJcO7tjNr918Mr59mKz
8uP7i9cB28B+Xd/s+svNpBYT4AR9i4q2sMAKYrcB1FBVzelckkzW2p+PsDFrmJFY
Rh+pm9vopC4brh1IhnbEO38hd1pP+9UvClNuR2arZyHXvYWRYM8mL3Hbjaqtygh8
0RVRzBu4LpVoWBb1fckcPdEKiObNV73gx5EAQMncygaPNd6msSI9b9I7wfS48tHx
GmE5ofL0wDLctqC9bdplxhZrSFkdd2ys89KQOqsLt3jFgfP6hi9yTW4WBYuVKACs
VmxlyIyAff0OJ/ohZ5IUZJ3XZhqYZFP6RwrQ3VKeCsKCToudNJKXVbx2L7EqB7KH
faAIChHb4ZkgzK/qT293BKdC585kcgV1cu35Q6yPiDnupskqHyIX1URcai4q+tPN
GmegwWELiZCZDwIKWjmVsTwVYK/2NCo1f7IUOnV2NTp+/3gCoWBe5FsJoqLTI5S/
kLMXX15s+Brx7c3woCXyEeISkqOJyWKZzXZbva1era3n79/bd+N/T6TV3bAyeGaB
RULy8hOsLQYFnkAVFUKOILRKT+X1EA8GvnM5Ne4/wwy4SmOzGQbsziPNmNNFU5Og
JCTheZET+mtWsAm49hAB52ETd1YiguuO0LyrbrL9ka2gEgAraQ0wcFTmjK1w0044
VlEcuLKTlzB8nGgxKvRs8w421Cm32AQTVidgramXztUxahbW7DdwJ9CTpfQVAHrP
OS5KvVPG8Sgyn064iRa9BJfMB2Sc66am3+QCJgTd2g/XWKMOlErgQ+rZy20WhKaY
g/Ahwa2syQfcBTCJOqxeQaziqHATlplwIS6GcfCBE/RBo2dVSoXVR6acJBV0Y7Ri
UWOY9vATu4JOah+QFK12nTq7DJ27Ej9RYoRudd5QUS3by6BHcSz3i51tIT5e10V7
Txie9OVm3cCAru7pN/tlFS1L/U7xnh3C9ERcD8lqv93Mo7g8NFtOh2PZGIrSo6rx
arUP3PR82JDie5cpTAHmWf9IvQivCoba4sX+7JnJGj2p8ns3wL5rGnXJvp0dV0jx
BNFMTQMxB+yPBfXiWvt6zrhFhtxI4JYylQs1Hh7Q4B5+FNl9KW1fX4nvgM30E87n
Va+A5ZvH/1o94aXKPi5ZZJL2xmp7ADFQLLEmHzmcMSUAE5dNsB3MMjT0ajcKucLJ
pbhHr5x5OHkPzaWpIy+U1DWOYqHq0v8IYmobHUzFvdstONVumRsanqBfBZpNnpoA
820Ez4aoxvica53FQU/S7KaamaNkyO+Rh49KlT2awiT3tnd3ZX39HuqmUUY4V2Xn
naa/nAIez2b5i5Sqq2gSXisD2/jgGGcfJRu+V3iC+EetvBVqYCv5oiAp0EFf/3gK
5UCj2xZvIAIgQmDWLxWTCk/7xdcw5cWG6Zsx2c1WSYSuXpwrZ1U6rC0Z8UQ9NaHu
BTfUR8Zw4VfrlRn2TpMJvaV0Q3ShXMCzWbmwvGaoO7SdmIZRB44nVsYxX6nZnrRS
MUbHCHw5rmm5CJFnMhOqDGFrrVsv0RjetKKDOpOOXEYQje4fJUliRfIFHeHWnh67
XBOTFnm3B3oXa2mWvIcKHS+TsXeScEeSAPs3ijHdPPTJCSI/9XGiTaKh/7B2tha/
js/eaOCh9XVrZKZ7frbt9iL09V2cXArcC4m+jL7Tzw2G2GlVKFlbZy1RsEKBAWJ9
QUTeaMow60DvjlEyFxjMOaQJHYgdCLbUY5BOwXm8/euAZad9wAyN+WQpbZDdvZGQ
tx68C0FYz7LtgBxVFBGeat3E1rV5ynu2P01OKZ7hpkwz0e9YHIBrqI6k8awDj5VR
4oVPO6U7BLbrTLr70eUYoZiUNkDw1oBtlYi0f5h1sBfaJ1R8PLwbKBM2WmZ0OBD2
uva9F0EG9xudIDOJA5Bz1ZGw0lccSFKA/TxWoaDXp0/fqsTpNsnuTR/GeXQUD/YI
A4HMiB4vpSF63XMP66hWAx0dh4KkostoXZfcMPWYk7XA/mUZTBEPl59X7CkLihnh
Y9MMQrFDZyQ1Tq2jT5Jp31dEuevAej0m8QF6DOr5ZUA/2P2feqRk+69WvM7MFmsP
SIxDLMjaeOMN/jBzWtToM8MqVUlO3R+/i6Q6lm2OrVnGBL1+cOOZX6z87l9U/9UI
n8vKHI9ukAZ2gdDWPIiJYoRzClNQXXHk2GHheTij9HLAEffDriYUj+Ra73VNIjUm
XwUUpBtZMmlvA1dVVK30T8a/XYzSFilsXsOyA4iY0cBnJvA+VakB4yWmu2QNP5p7
NtFTHKLoUedatUqbxf70V2pkp8g3y848gntI/a6n2Odgd0yOrazVfpXH8sDuEkJ5
IFJkWoZqJeBgfSArc4lLiuxKF8+sf2Vg+HMG7Men9VcAzLR/inFhuFZIGR0Ex0Wb
WYwMR+gTfjYulsMcWaPtHas6wqlJ9R0jRYrO4W3sD8aEYRi63i6S2MsS24vlSukL
As3W4WArUE4HUubj8mLIpww4d3cXHBhEt+oEaUGXl3R5zaOf3r0HMB0FbI7EaQQG
PR7OsCm5QaAjwVKnuDfBUvs1ykVJhicDZ+z4dq7HHTJODahivEN19aZZeJiEzXH2
ulowQ8LfXFKeTYqM2e3gpr5xE0oGpQ3AMnhbktGRd1IE5u3my2wWs3/MoUbcUIm8
Z1FeUyTFIsFhqC8YNunRBkL+alVPnn6I9PZld5HiXMHcTKqHUeZrj2f2P+BgEBJW
vLAypbY3NL2LcWk1z4gGvpNXyTQ4hy6HHxyKDLfPH+Gxqbjj/awNUkWHHasq2+yp
zteqU67T4bgCThuU6WtzU9nyLxik6SVuDeOw4hd8oK79qPMzUybvlinN/3qnArQM
Ih5OpX0zDgtImEJGYEHqvH2+uvbUohbBAn0yRF+Cpsh/R5bo0Q5BSZDCDdYUzLMI
5yQYC8P6VJ7/o81yRVpMyhNP/Xv1gfIT9iXFWoU6uoJ4WUdmW2fDwnsv1Q4knmZg
D6rA1RSF0dBO9QzC5m05hNScEi98BXlzOqOY4o8arm1XkZIvjUDjQUao7UZPMEOh
KhAp71SuJh/hOkE8H7znzi2MjIGiwYzhKqcdKVfv4dHkOHcVM4JTxVeHElbGCvus
2AMSnZbFIWg+7cgYygQGUVkgCj6pPiFn2beQMjO2v0ZaRHnebaKWJtSKYvqOx7d9
HJ5ieZ3H7QBJEem6BWY+mQrT0mqn7JdIkKUTmHKauMy7xJ8Xu14CKcSuYNi/vs0c
O3NP5ZuPaiqougqcKDwukk9osQOWmGE2EB5pyULa6AMDaqHxVCsQsFz9dpAAEveC
PYcQ5QZzd2u30mtWQn2IOHYOzpWmV1Ie6e9e9a66yQBNoaQktS08sNw9hjWo5png
PYZfX0Aye6qP44ob4GMrRtPJR01PmrupQx4twV2OBxewGsIr+F7Z0Nk8C6vubIs5
fd5nigCp5GhIQ/EryvAzoxqJXm6BBgElNw/iyzXojkJV7mANAItL02rUi5GFhlk7
5Xz8RaYjyL5HE/EQ8KjbNCtZBejjueNXcr4XXrOGuHfhUFt5z7OZfBExDsHrJO+9
kRHhgjWoa121gyDIK6SuP+wd0gRiZV7LA+wkNqSndlQDriTEO3XAQCsqlGdNVWxH
JH67tfATiItr+4xoQ0fhG0BwlumxwlULT6i6jWiiVu5vVmmJ3p0ynYFDVzjBCyky
pwDzwluSYR1h7Ip/nXqB48R6lBYeLMCLoy/4n9x3zF4mH8xBNWLJa8Y8WllAiWb8
e4zV1ho7CmUpcE+9L2OhBmFKaCsWTm7MfFadgVjwC4IxY5/Rz7ciKR1o6bt+OxZ1
4wEwTBIZnea3mxXlQv3Ox0IDCMY7RoQN3/TSzKb4vkUBwbkx3VjdCBfq1f6ZCg8V
KvTkGvm+2BqJKennzR5botwvNiYjTYf3607LcpfmxNi5NdpQBGuOHkhpu6OWpL12
/uoFKqxDa2W6vqcSBCCmuXkdjgiuMt32lpHG/s893ru9gGx2j+btnsNorsA/J5zW
mTDLDtcOBqKAJBWDWRVpiUNOBf58YHc2w8xUgyQZDQ/0nRWXt/uTHJA838ld8m+N
`protect END_PROTECTED
