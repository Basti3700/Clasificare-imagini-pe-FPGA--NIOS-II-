`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/awslKFwaK3PmHJn4PDAEPuS/QxAeWoABLwMovqqEf10i43t/JtnG1dcTaaaZv3r
eW3QZEWGoZjFUrx865Tl7zsr8FRbbF07wPdVhx5kw3NY81e9Iei0SauH3OSG12Lu
+vqg3kDafvDgPPaMb1Oz4KBbmEsOWGmWQ1iIoCYuZ+2okYeA0mRstSnzWt2lmK7h
lMJFw+wjFvMOUcwuXj2qf2qArt/2vFIjSwWdjo0C9Fj2uPo8dpQi1jnNjSDWJozA
/MG+0pGxp9tfBypRTx7M6C1HgWmjQqsbGKnpy6hZWVGDN1AlCbubRm7QKfkvquTr
YUfT2AbuUJF398WLnPBatTEhHenO8pdqemzUqdguga9VbSjKnKhVjSqNVJAK9nNx
Rh6fFXRofHKI6f847gsnYbJQbv6VBT4gelquDNKJ3rowcdL1xaq+2mSC5Pt+jyBh
eS7aozMduWib/DCgxSiipzHmUmDkhjd2RhnmHdFtiBWjC/byqDpxKM52LWc/FBvF
0hmUQoq7mmKrEar5BmtbmNafetllT9uzWBUsNtJ1zrSQ3yFSv9b6L5RP78FGxPKm
Zpm9UZfMmdV+LItFwX9WRTm1/xXuPwNaFlAfb/saF19bfEHJe/XHxrGZ7//SdpwG
GROZeWLYckOnaqhoxYcujmOhZJtimFfwvBTKyaNo8oZvfA/dJNwFEFCQSqcvN/yO
EyhMrCJAiV/qQ43/KgnZyI3FcMy/d38iLPuTWB5kDJtqoN7EFasY2znglaPkPVnW
eWrhSMGIbU7z7m4x4fzsFPQ66LvN3H7jE1gJH9fBu4nxFmMoMaUMnP5ioUsBsWY4
KRan5FFvoBrJ7/kKGfZPU7PJNv6eqnaqzJKoN4JEz6QobMlf359pfSz864Mq5BS5
FVWwmeCcB6JdSMWcKag+zKTbp9z8TXQlY6JzToRaAiMwbdTPqc2gIyp/VsoqLtcT
J6LCUpI82Sbx1JiviLunASfmrORlTx7pDiKFBnFfjtbV6ZSuJ+wbbQamD/9/Cpk+
IGJ4uTIm/KNVDqPvLJ+yTTlSP38Oda8PqOa9JR8HakJxrsz/IzvrOuHH5rihppa0
IXUlYuYGhTMz7ViukNrlMT1VcbscDlKFGxLLSL0ABPlqLjtdEH63ib2owU2/kreZ
svT4uzigGpBq7sGA2klZj7pzptRYJvBsqhjKdK+WZx8Cq+8qrW1zyx4+jlE4fWnT
xl6Wviy8rxPm4j/XfLbJ2u8pB0wIAkvYROE6ZBvkrU8mVVoWMll4u7zx9nlCfdN9
Sl3UFcAEvFQ6YVc06BSuFD5iBdM8nN8qDUSE1pT6b8YjyTubZt4kx4dhK8R5TFwp
4sHbeZLVsUG8d5BRnRYgd4xGrrsqhJ+SnBBrejVMnuzBN3IWS4kQ9wQR30296Tv3
IfymXbNdjy5R6wu8vMT485bIiYTfjpo+D6U09FJZkRRCThp6vp5Ot7eDvrWPf6ct
xOIFHcovSobgNhgv/wBcP6RIAweXt13Nj6SE8E10gjgkWFj/sj49oyeV2f5sG4GP
oyPfcy2YoC9rlCUEp/ve55RNFuNvnbmFvxrtqDZy8pC4bqcPbYdR1ALxaPocAY7y
J1Y7ef7FPSObf3BFPb3/I62uMhygRJemnzBIHC96LilYX/g0OWX+rgZg8bh9mlYW
exhv2CtaZ2XvvOWJ53+YxASwjE42xjmwhipno0WaoaDnuQpgBflI3RcWY11TK92I
1Pshkk4fYzPNDgU6gNy8EMNwVz7C0/rA68alVoXQ2E6OMQL75oNRlQLAx66LR3uv
LtngkVUvNpYufebObkVGhrPdiypjXGFLTjGp84O46BX5IRKykMtE5uoh1yqwU1w4
ZDj1T2OTrp8UsUJeW5HimkZ3Ja1bXSr1/FJ2grlSCTOJhENpgrpcMMlXQF8Rwa7s
yJzmW7FHZtNhDdfvLnsA7/hLBiIQitHPyiGUztRaVh9DfLwfJY7jABzYxF7q92PM
7jY2O1G8y5ZbD5PtZbygY3zcutAo73G1Z9jHIWWg9gPSrw3cE0U6opRiRdgWncrC
t3iKPcURNIGLchpwDBGWF7bsHBc/xeQ+IRSVujddLZc/udCf7ZeVBBtZbv93B3FR
gFFpyjq930VsFHAr112WoE+A8S688wMgEeYqomfwra6TSGYNUk5HHDH/Zq/wt9NK
TsMOKsdLNqw1n6HVzr7mKe+MgFwhyB2dossHHvMG0mUkeaCqarlBZX2PNB10Q1eA
QKRnBnjwYwB5RQzapdGwnAaYB9K+vpzxHkVjwbXY09NRvqOup+yi7/3jn4gvEoUC
a1Sk3EGyOSTM1yjXlN6BhPdq8vYvTeqQwK/HS21PkIrNR1MwWiwlHd7Lr8rjoQN3
cxoW2LA6yMrH8YytG0T49GKZH3RPp9DWqxbYdPlhiKyx9zKf+Wx/js/42aL9ohKK
Kktmv6UanIBzp9wsMVCXqDi59Jx2BA7rf3huym/wQ04EuvUppv4gAN141w8KDOvw
5o01OmyWcYBxfaNNMqry6+SUX2g4u/dKsg1bZoeHYCHWGla8Gbnn8ZAulOEIyhVa
sEoCl9c/IiDXfqAE/QvZygYjrtIOvKcLQXq5G4DHrrNZS8YAjMG05SB9gw6djwbM
BcmVtiOWpICcnqkCGXImWF9WQCm4VhEUvzI4hwzIUlZCuPrh+dwIoQaKk3v6mcMX
RNNZnMpHQwPhYOYCkLWIPXNMX43/CgrNTXWGfhuL3F4gQsVWGDmuQ5+6eu041wQm
nQAZ28vfkkNVk6hjqg9UjOoVndFYDn1PfLAuB5WYjLO00aqiV6WgVsJb7UrNnEGX
r0yxr2bM9oBDhq6yQsYCo+QywEaigwXed+yJFWzoTbkqExkYT0S/cM5npyQrAYXi
WbQlLTEcE9tuD1tHpsmVzQc28F1o3As5eRBQ0Yt3dybBZ1QoYL59kilX/ADzmZZ+
CEYY86uSLfMZ3xDSWUZ/q4uFanutND0Ks67HPmef0bfZdmhKhrQT2AZ24F2uiLGc
OheYyFXtIgBKl0w6T+XqjbxbP5mR8qncYFfOSZCewQscajl/WLMrUVkBNL2crzwt
tSPkktuYZNZT4eVjbk6z8zEhmxN9js8cjti5rTnf+6dw6j8JeZQkNJe/4nThoKw2
Q8zgtiIiUaGEoQYtJSCIUurUsb8BuxT3PGbeBpWxIQoU4Hz3gn0o2CoqgE1wY83A
ZXDYdL42rIkAAAboloTA5BEHG9pqbFcb096URPKEx3MpltRAPoqeF3O2vbfwgNvb
/sC2ICY0jIsTMZbFgrPj8ciueNvpEu38qHJsaVZyA7DLqNGiSAlvHZ1z8oKOKmxY
YBasYbf6+PxBYp3BXdoCeR8kkif0SFG31as1btmLfoVZsaBXOVtP24mT28HQu/GB
9ixxfYblX3bxxPRnGzDhPe7pU/Mw5toOdbPkgHljn9DBA9C8r0iKUGDu4Hs8wFkk
FqCw6bbbEaJHDVM9hOZ5eob6y9c6vyysIkmvK4xpZaIoCNxHjrjshjIWB9XSA9hC
g8KQiMkMAaKdpPJ0MW/yc8lQTZr+nfBYA8Z/+nZCts1s/oIBeZJhd59k21kDMbo4
wkCoGrsmwLH7ePopGiQv1UTisO7dN32s5n+SPvFQ6Rn9jxvTBxHdsQcTXhZW8Gdo
GEd5YJaTZXVf1oY7KFr0UK0P3hG9PleJ6NlUGbRUDAZ6q0/o5KXV41pm0D/sKXBA
nOEaM1sArVRQ20tDyQG7S1ik/rIgE+hdwBEOHFs/It2viwkbYnWJi3njYoCoRzcT
0SaYa/pE97CIiHBuccHXELlJBWjbA6/7Lv5HnZVGeTcM9H8WIR7dKCutvdaG9MyC
VaG9Kh+Th3ai0cWLxSKyhnt6wrrxLy9LVlm6Xur9OK9Me/4goJePMxFOrPhHaeR7
DIjRrkYK2jv644k2OJZaTMhLhN8my2tNMC0IDJ0yCk+SO/vF0VjbB4P98vd8zjaJ
gvfSfgIbjDiAwwbJDMXVdDv9pRRjC6KHQIQ7X8/qAVTeCSz9Ich6fUHNho+I4dOl
mkxPOOd+raul7cK6UCKVa4J/u2+wZSxZeYvZZ/542+8lCCPHTm7IycwLXg1AdI/B
Ry/uohE0yvGHOBq1C+vjjBDGcGQdIE3gB/P0Z40PzWjhpCAClyWnMBcrGvG+vs1f
wxG5pmEO5Tm3w8mnK2Y9DCUwp/DZQ89dvMg4gNjrWBrdKQXtNHZt9h6FYOU+SLjc
ezCTgxuPWXbn2MHHPijjAAXRuZ5jpj/pO8kn6SU7bGMdCnUJujixktS2fOjC8muc
5noh3Q/UkFrlVX5U/A5qwPlqcnorhUEFgkEoRqpKBDdSDOr9g2/TUclRodpgErWi
p9LIwUJH7SDgSZk/AgMT33VYpR1zb1jfBYXO6jLUfvw0WVbmzQOaURK+LVwIhVrD
z84hNx83rIkLGM6QwqrftQOR/omkzTJFLas+YMGE57sIAc5wkyWZ9dV96uQpkB2e
IxfFW/M+gWQ3J4PUutzxVsWF/PJntpKqoE2rUEwnLPN+DjSrwuB8C9pbgFNhr4V/
Qn0Te+HIcO+BTEhOHqUwfHcCvb+pYkacqbKqJH6rPYNSRwVD5JIypLBvQTZJHHdC
rcjXeFTx47HPBM8u0jLDXh3imCW9e2i1idkmpZO6ysJomFvhnCpkZYOXadFpbLHH
CcxemKyyxtl3PmH2MpIVLvj2x+WfBiYfVg5P8IY/FZWc4xjFm8YObVOmlo8DPSoM
Dva32SMoIeGD/SY48k2fM9/2nIq/XeHl+Xf6q40QGTTaD7xKXfmwVTwrUFYaxhuE
W7TCNOdoXBaRjTGpUcU2i6Am7XJ1q5ABCsbEAcUWPRlXDidJSZX1X+esTkVUUU+2
4N5JUR4W2aYUiPmMpZzozFdHhOBF57Z+DS8iZg3o90+PkXw6T7oHGtrDAqhawRMm
9hGlQc25S5TXZvDSWWscaf1+XBs1E3bnD2bmxBiTgpyn4+PVZkvusiNj42X+BD4R
UCH5qMNqaFDF1oc5qeTobPDufHeNxQxFXZIaZ+LSwHpMFBxaN7OB5FGoY1RIVpZF
2t2QRNkLl+XVaSVVqxzCGSyjznPFy3i+MP5I8w0lVvu9Rs29+wFwzXM++8zsMIsd
j9AiCKBOkpy/Dis3YL0NuX/JwYZvH/eetBLAEGwIqfdiv1UAYekBL+Yfqp8tjMiH
/0DWgTLzaa8F5juk9RSZkWQwdSUle/UTrS1UDQ0slET7S9POTl87ZoGgaeN4PJOx
FgavhXZqqyDZWYXVKA34OAp8Ox78X7/uEWUZZ5r2pZQzVFgEKuEJnBD9VVlYF4JB
IUFk3v4k3HDb7QdK7BQf1o0p0Xv8dsH2J1bomolhThX4CmELRKjX5L4NRLWEPawG
9wILGb28x8OL6ZUmn37EurxvhwmYrSJ1RAs85uGq39h0SD8Dk47psROyLyxEqMhD
xEXsD/BRHDH3ZX97ax+nBB26KIbRpnu16JwBKWGA5vr3CtnigBAzG9nEc1y/d16i
m6GkeErIOSzgKy4IUc+fHRmvbX0u7EmakXBBnLFTYMqSA8wYB1xhDruNvLDlfINx
vbwR0n9YVHzMmzBljZnxrDaLamYaGqTpAB3eE9cE5WFP3FPwzplsBHCWy3KQlvjD
eJGvJ8PrfJVOR9+dE/UBWeJ48rmTN7i7dl5U/8Q8TA7ZtdYAfoEFVif772WB77vE
ahPEC95TFepMv52a65VhG/EOxBP73raSh3vfkPfVR0EGxQbdNXSU5duojJhXjSko
NW2d8+T40jPXD7K2v1/gs6Dy1tkC+7HJCWklDFmCgD9thL5FGO+OCjdZGR3X8p99
OBZwexsp0PYLjfT20VzquzYDdzmGr/+BNgE4+Qpqq/Y1Si6pb3PiQmhaNFO9BlYJ
vjwOOCz3ug0GO3l+VuIBH+AzvuGl/OftUtK4q6q/+CdJVrZ2p2IPdGJdi5NHsvw8
H6XXoJrrpOD07E5aZgA+zShItNwjiIIVymE58PEoJw1knUdVP2zZo4pi4rwKXNPZ
Y3JgqqKqSc4/IHoed8WJnwYg6hKZBtUyTUZRSZ0OC7ZAoKwpBbHjTtzTv/P3yEwK
1R4fivau31CpoP1wTJPqv7SOIlkCcyyxd8KpKDEG9NiFVpC5g0CZUP7Zm+qBqgNc
4uGQUIT9vqxsx2kdbqFCLbjc8u4UJNf13ql31F0yFIT+otQ7KgvtUAlwjs/q9UxZ
zOZnZPRTuJYwkPP0sjxTYai5y6vlttGrp+JA3QA5zW28rH9AjUtE6No5etrkd2I4
GGNN5+zW4mw+1kkQPGG74n9+KBsah7PkML7CDdXzhA+2Ucksk6sqCEW2VNp40BpU
2bkg/qcuv49dka9CyA1xD4XbLxeTuxamz0NQdxiGYLWpaXmfjJr9pgFSF40W3EPT
PKcxmhtHifZpSxOfUTvVq4xFIZy1mew2TjQJ+T5xlmMqL1il1u3fu8K0fHJ4fS4O
6oH5BirILIrBzqlYVp6bBkOgWhH7O5lMQ2DnY8E1452SPw2pD6UK197fOkO9r6Y2
7K8EMDhIANyEKcnf84uM7W4SVr/Bn4soeBRoOR9zdlGdnbFQSFkm1asQJ/XlLkfP
n3lqEFC7pp/Uz5oN1Pkl5qlkztO8pUIciHKFBHVSBBJnU9AmGRxYos5aI8d0rYKG
A3aA+qkd0u1jyfMVz4MiX+XLUql/344jDQEJE3ak0Vb+/78NQo+F43piWNClTeSC
PkSqdHy6o+TGvJITs8sMgaKTk0DXDY8/xndkeqPWrEcgF2U58wzg5GV03O3OX/5S
wZ9yMw1mLhcjwyHhKs1ycPRyWY6NVQtWXj//2uTbAv51l8DuBcePHg17qUDAu8h8
VBQiiwj9bYVurb43yWh8bfx4WvWNl7ZBIDs7d1tcyTqQGmYs/fmecgcuHp8N7Blv
F3FT/VrmBx03V9l0YNF+GdZj3QoN9fBufs+HeAiZmJ3ClUqJf6l2lW8o8H8ely/U
GVyYGbYEx/GUMF+EAvwsVjUnQiiFjRdJT0FK46HPsein/a57VLd9hWAIALuCUdI1
Fi+/q6zpu9JJHmqe5HfqNNo94HWx9wNoHvLN5Z3jicGGwZstJn+aLciDomfSLW4E
6P3pPTn+rolSLZASr3ZaymU5LWS+p4HVWRBEzJtbU3nMXyQ1oAyPL0/zYD/+usso
KjsFIdGF4IlArnDNHd7kdrs47EREc85GbB467FfyRjKIaulwg8T69cTDYzn5+TiI
nj3xRKz/+1JzcxpjuPrX1RjxAI3YIBYqFUZfQ4i2KShpomQL/0u92UMKlieeyjQJ
Z7BK719pjt/WsuzYAA9998m7J8gFCIrFQWbWZDtWAancu+jUMKLJ90CM7/qwF8yT
uxDhUemPkaHAvgOwlUGGZ1qXclRSq6omJse1nPr692YEcTcRUEYJDsub9oX5esoP
0ixlIviSvmCRyi6fQaMFNSdIO5Hg/vwU3d/ZNQLxLd9ibUIBELTrKMeMUxVa1rIu
VfkbLwJQcthUNF6MysLbsmx1KjZrvDoTN+YK+mRXrWDtJv/hT3QQIfgriY7goiZg
hFuqHRQI2gHnXOHWA4bp6/BAIMl68MJxjQ0eq86fPURr5Ydv4jqErbEG+R2ON040
QLw4lfIJa70+Vj8YWkvMqGWewFbVyVk3WCdC+Uaq9JzyoktM5B7k4rMDPQlV1JRf
pAzQxl5nKY+tVNYXGh3Qpp+EFrK+FX7jH33llnVXESFi7BLTLCzK0yRmzIpqF5YE
XmKIy+L6truMq5l8HxTBe6S9pE4Fn8ZRuBmnIWrdyJvET4xmujyOHiJmbAALZlP2
voqJV0dyFY1NSytH9I5726sgcHcYa0sxafNV5iW7CRmwXBmULDqTusyJVvlhy3V7
BzemzjRafYthI68bhsPNIWR1aGU3qUemhXesBZztso4Y1oFGuowSwkkBSrmdbX1Z
G86+TA4UWwYq/IgbZ4B8Sflb2UTUmQ9m47yQeEGMoh6+B8sODewb4Fw/Y50+kouX
qY+u3it3S3ZVfpty9cr7wS/WoarIEucRV0fUupIdR6ua3q+1+os3suSSn3fyMmrO
aU6txs6p6x8AnvZaU85/X2eA/Hx/XoLmmJIOSsP0f1kQLCon4oLmSlGLmf2eNDdi
35c/rz/GBnZ9+iE2ZpfaVSD1fiMoM9wP9uznfcaxMDb/1nx/To4hM8o36EKeJs7Z
zY86ROMaoPNJ5HXwcLjoTsx5ydvfzVSRnJZwYZ0WokNrJZcrlqLyZpPlBy2C9HoT
nXYRnkG0YUNwsrqddm5+awvFKCx0JnvgfT8NRVOy+yNjRcYQtYcobIRLXAwDYUlF
g5vWcKcstbsJ3EkRq8FRnhYZ/bMsGV9CPgJ6Umtv6Jq6WqBmbuRVvsH6W5lIu17l
TTtfVjdHFvPPuMRtb6UkxjdFJ3boIJ/3j8b9utglzGsZO8sVsFCNoCgia7q1s0uN
PUPgVrURi4OHQNYBbh7jMpX5TUFX41l+cGnDgzvwWRbvugwWe3ifPST7GlgAgcZW
/2ZMqdy6wqH00pWni2YXwImn8fsqBd/Pk0FYYCw10/mGHK/7438Wz28u4JCrK3e3
OS4dl4ZSc+X48I9GQhptCKFUJfHQ8HIzNf66HdKOap61qE1/5oZQxwjmwZB9X90o
43kjwKRlqXvadQALOFAUCjuPNTxeJVpQiBdp+AKw9bx2xD7orT8UbTmFTxBSsbhT
ganf4gB+aCHkInYx0Z5pcpGlgoV/HHwlZCY9lLB0jBNQuRYAlqaNXwCed4DlG5xF
AbbElWoTGDGUkx0WBevBaA4SSRHRV8QkSZaNeKOQyPLJJhUoxMMfOjIBvPo6WYOA
IvbWAQFSSV+RK1N7kyARhMbZPti4ZBevFBJhs9R6nRPkI0NXTDMH8PaW+/Di0k1Q
w4MeqMjm1V7kFaCJTUcIZt7CK+aOi+0uM8ABn1g5+haEq/z4K5uPg+eGLS0xdVwA
mtDU68F48ha3AcrdHuLs2EjaiDRb4FO680wJ/oBVS2E6QVZ4xdK+5mScN7EppF4S
ZZrh1hsFOQfp4E3NY7J82QACkzbXkJedFcwe3FDKz7Th1rBP2osU03nOtr98kUVM
QmLM+A+B72DfKT48dX/CjHUUgEhE6Yg+aH+JWeMqWx7EiTqYKya6+7jKZr3x/G/3
BuWliEs+hePcpP+2elX7b37ZlJNDYGe1gUEMls0so24ktTN0pEiq90W7DDaB5Is/
SIOOAwzctNMPin30uXSdfX4SG4EfKqoxfzoGgCLWKCRJlmKfO3zFiHSJ/jf0db0k
TThxQsqS1w3pCXY4JpyQ8oRUdlD/Mfy7o9dbCqWxdSFTAhmPL7YlF01ya0qf0iqE
VJoEu4G9ntgznJyyY+htRjsoXNJkRQSW5d6j8kFZb11ORhw+dG4MU/2gqfgPyHoy
b+GKWkvuGydLz3SLnKZ1pKd565z1B5slDmLZ3SiXvsoo5tsuPcBktbJgSRJNmJCA
NFSxaF/0UuUJvrWPRtfFdsAJQGbqBmJLUioQULMG6o9wW/BcBYS+tTe2qrU+4IxK
K5FVkJX8SbS1mQnhBYXt0OPjC/5wyy53rPYgRwZ6Rscl0wSE+061HP20zyynje1B
lr86wChQX/n/jIxx0EzZzdq5jufFUJILNzzk0p4GFEhoiriHWHLDfTlGpXPJCWJg
bXJlg+37AkXL3jtaXi0kBIXOMoqgLqT+Mkad+0J6jvDtp2bb7kDQWJrLFn7YIw4x
Q+H/QOnNnsBe2lhTD5s0gVzGRMdaREANECTKoiykTc5/W10pPIf6NOtGJaqAVe3i
t5klvZC+zDE9Wx7OHPqicc+xfMCDsFZvdjwruAIDQHome7efxrF877UREOCL+y5A
KNyZ2djxTFCHp8Yt+ubJd3bZr1XZ7S6Erl0ahaGpOlluht3lq2H1N9tIDXRWtgEf
aIjwCq+PGbXQhPfNr9SOXV7hZwbtdVf7SHuL9rFDCmEQ6pA9/AEJ5648zWx9lEO5
ZjwBDmVEIgRNzvw0vp1Lcq71gwaxo5f772g3gydrgqm05a3q++4kmCS+zO4rgXTg
aUVk3SXRV2TT+qwE+wmKn/O7T5bcWWddxwhi1eOoBM5Kg7g5kJmAPHP2Rh7wyOrh
uHRlWBjT/Bev8ecREi55VE6kJO1XMdmNd84YEneyJZOUACMk4RMLrB8OtX0pK3FM
LcGOm75G7MLoxoyO6nqlsfri86No+cXRgrWLh8/X72NCtuUJCMhutspgQvx4h8tG
JvZNsUzbBW4xQrXbTHkyhkk83k9TCLRLsWqLpzcNE8NYuCLfTTxtpYNXCuUcC4Z4
/ZD0ge4dE1VxfW8grB2pf6vk6GmVaDN0/eXb9ONtmnWcJ/BE1C/5vOD5pznYh6/Y
tjvopWNMwsNJTviat3K06huPxJrHRZ8Tl9CkTK8Ahz+PMeS1W82NgyMXkKyghBku
Mp5mGvCg4tYywa2rnF+2rGRSgc3okODom60nTwSqeacXTvt2pIUtsRE/ajbbIJWb
WC0KxmB86SzDBKfzsZjWeYlH/KJBorWBwI7HaNh4GMfa3NtbMT3i9F/mj5ZFPSvD
UMP4oKHkOb553CsY800NlYHaTpQMK+2i5jf4CpCGr0VRWN2wMVKNCHi6sAdvwnE2
9fNxak7zuc+HHiP9e5oVRptQ99u3xJ/jtdVh8TKeOLh6Qs3yAvJvQErEzvka6fLp
UKgQw8g0Mj/aVSGy7XOBv3MeOZvDGGHpetfOMDeUTNx3C+odY+SdNMTGqemdsrw8
BPmbgQIPK0zbn8JxTTnOJbWNoES7ba0S3tD4LhBKQguNzAnYA/XFhVo9503Us71E
KrUz/RbTKKTi8VjGpNeWtom59BIikzqE6sBW9xhv7+Rotjhmxg5q2aEJs1yAZWo3
mWCnaIRooSedCF7pCUHQaJFycvLVV+8NGmR2pBjIyrNb1aT4cGTMaZmhecxG9uur
vsec3O9jPW9rq+CDBqI/bu8C9I8HRZubD2ahahfGrbZws8SSBVg2B+51t9qXDU6F
Jr60Dp/kaTnG5/W9oG1//kfGbJ/x2sFDKRHX2LSzAPtYH9ClnRvL26NRZFmZUUgV
HiGBP3VW76LMugkRL63Hl0oY7uPGZ7wy+OTw/6/RQtstel5sW6Qkqo6zc3AhFdPQ
vqHSkeY+j+aEkWOiec8faVyWAUSyHp0E25Gmf/XVjMlUijDBoIoon0rn5algxDQY
ZiuUVX3uZKEYmrSPMFit6qPzh4K63UJzJu17XDl5WsEEnhuks+4uv+oHlr2I0QS0
NRr49621XQ8u+NIBVaJpMb32QXiP7/9fGlIZB658tz01blRIcxftZFgpRobFem5E
dV3t8j5k5hdjEYoGoNJu8/jiPCCM6g5fPTDBw81YqwqldEGUQqG8ywyAq8DU8xbU
9viW4UNL2jXyIc/yplpIIbnkUY7lPJTh2NCzGFBnWdbTXAcJ2V+q2Ay6ui/AFPXV
LjvEjZxBtv+W8zm75xg2hDZY77N7y86onNsot4VW5icrDBfaAMvOp2UUbCXrkoli
iv/Xe2+JJsx9RLtLtWJVSchfG7irKglaLethd6Memsc5EEZbMnFoL6G1r5pY6LO5
uocJCDZqdn8r6QezFCw3GiLLYB3j5rF8mcyfYq9L5imECP5quufv5tQyRyaoiyGC
/ip8jeFAcTvffJTnoK5i+EiIqbSXdmoGPolY6GnqsIa9fGhn9th6y+NdhMX1Z9yb
SWiF0b0hC0oFzXS42urIMlFBnYHuNFBGyvWfq10HF/fV6ER4ipLNBok+Ax4THrt1
s3uFp2dhpzGbRGkpHEigVTJThhP7IblEbEXM2Zg8Skg/lO20GNsTITDRFu7y8HN9
iK5Gm3AvhG0m+qY6VnQ7a1RcuRKv8cwoWQoq5Hiz8nh/XAMtimTV3A2+shpdHpSx
n8Xy3MOQ2n1RYAAgoWjjKtPc+ALd++C4FH3/NPvgVJ7g0hTmWHGwETZj4f/ba6IS
ynZpobZ/LPbI1COhofXO41B07+S8kRNL3D1hJQGWVy/xXbg2Rhap0UQ6EJAIXNVB
G+90sUGpwzpvGYY1eW0vSO/DiEM6Zj3EWOJ4DJ13zBStTR77f8O+tHe+0F/7QENA
`protect END_PROTECTED
