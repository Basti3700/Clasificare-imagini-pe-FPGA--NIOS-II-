`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oVrEnoJ8d8qRn0+6gmuFx2pE/YCD7m91iZXgfN3kQcyMKzlClggb07alDST5JHTA
VtCP2H5BrRK+BHBkByLICu8RpbRuXK4qkSvwntsNBISRaiIlBWmUeN3G6/umEb66
/4fw9GbuPA9h0T7fRUE3jlYlNIClrwmBpstprdpuvpxIU+REphJJQxO0YZb3cP1n
ce+8ZMiN8pye7NZpD91Go/B7JH6CKBE0NIoIGSUEFHvGz6q8XrhcXOvShpwbx43l
RqeYoj74tvfwr1i0F1F9CdXyw9vOER6aQwsG1dpmZYSbs1fMuDr8T54xbJwAznif
JFaY4rOJ9iTDK/2ZkkgN76QCxUsfbjYv6PwB0NGGjPlUQJbdRD4/d5Fvy+BKpm5C
ZBd0OhCJAWNCsb72Sj4EoH1mieneYZLlgCYgKL4NvRcZTJUMdW5k4yUcNr0HJK7j
QoCp5DumVRsJ/72Tdeq2bFY0moqMvQj/E0lR7f9ay+zho/5nnOjAs/V69RbQB/Lm
`protect END_PROTECTED
