`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dCBWl0DDMMWWNtjfwWArAjVXuWSgrkMbjreBTY6CxbpBW71tVMj7Pe20xd/xVTxd
Eo+HYWvWJant0SOqcz/ZVGhNV9Zo4/szMjFrrJbVIQueJwG7WFZnkRw4fevVIr17
rifm/moZo1RFKyGCP3uz73zvdzv6rFOQZCjZl5gc7nXxmbNbuk6idXRqLnlQmBmo
Q38lzd1ETFyWjo5qNNhQT2kfKyVOxYR/QSYBVRYv/wE=
`protect END_PROTECTED
