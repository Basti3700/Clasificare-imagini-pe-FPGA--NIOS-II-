`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CNSK6UJUp41Ck/j9tUx+Mnu+YvreM5jiXwQFiePG5fJdDn180OSiTdG0l6aoLHEZ
uj/mpAHojTnPEGswbH18NFLYU/4gsIDZSlWdtaQFvVdgJIHuPjpwlCryeJc5v1Gb
tZbigntR8AOEFx/MOFPyMMXf6mnzp9oiUYw44V2o7lPOKbROy3I8yUzjl4raBECR
1Jd98cXnDtpz08JLjVrMbo4mtDnL9IK/HzpJDg9mbYTTSlnMaCTvAEie/0k2l9//
Xq+KavB7iswqRxe/jnWcHkLyO0qEFJcNnhvJZ7S5vIlfay39LBUHMTPVhRDpM0sn
X9yoyQHV3J4Q6bxkiQ3oUMhVcHhdeaRiJEj1u8hyUcpe7Ut/MzQBbQgiMRyuhEtR
SAaD+RWhsnZJ52bl+neU3/ieuS4IODzXAcOQpSk7Wwvus+a2Vd+Nc50ktOCMPLKk
ZjpCxX68X3BECwgf5AYcIWdLBtezl8MDnffc2wrdG/pE/xY0oqOtsNcgQKL5UnkN
l1rnZPWNKTQZlrAUHjgW//6a6m7I9HHu8eFTZxqQ6A7jdE1am+VCncoTn2MAJvsz
ow+mCyfVRNQxR07zur8PMG3ef6gJLKw16PFDvtH9UCToaA4ORku1DdxwOM82PaZk
aJOlmHwGbAArF0oMEADlVRos2xxCHYpjIm29X8PbsadHquP5QJL3Dore4otqpbmb
7NZpmPIDtZ1if6AYCkDOaGVxQNQbuPtNEy+q2onCHeqzwkL+Z4uyvR7UCJMgEaZK
lCnYRG22WjzItvSkFOM+b9X8spXZb/sZOCbk3ytTarURoaUfIgn9Mn4TGRmBCNgo
0dul9VHx2vueF3yR7FqlnhFjkAJALDtVbk3IsSAo0UszVyzQGNL6jYqVVGb4lTY7
Ah5cFAN09CrhHHepq6wwyfF5oLGFpt/3JZ7oVyQvIsSSZR7OIDjG+GlgBD8J/fkV
kJTVnHAsfQIIY644e5sbnjpBn51iXCcsEMH6KjppX/HE/YIWEcBi8pcuen3TmcAy
oRdt8iL+el1YoAE9zgtHAQRDzVBDA8Ulc6IjZmEAWtkzf2nn4Y6pGcOOROXq0UC9
E+FY4ZWA+4nCprhCk+U/7xeRdcaX0d0PPDc4TGBKFapycbm+/opE2iH/Gt+ql6Jo
JlcKT7CED+Zl6ksbgaCSNIve7reMprffREhBkTItI/5FMYncLRMYEhXIrjfLnEr+
t5E5TR4Af2Ey9cFSG4idok40dM6nmXkB0La76Xef8XQ=
`protect END_PROTECTED
