`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6qUtYbYPT9RWeAoEz4NHZYbrG7r/aTCMcigSmjd6N0N+2Y5AUfzinJuN9nu+4F5
w5+9S3pViTOmo1a4zyv1MGWBfV0UuBmRFVJdwfZC9yNEHxW2XS73ececDVeYEuFH
/97IC7xQZ05QAFHKnzCIyyXw1eRIbP04G6TeEEvOn6tLOtDdPdr0AlEgWUcVzhzt
`protect END_PROTECTED
