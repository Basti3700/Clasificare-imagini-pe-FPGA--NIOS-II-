`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ksyyPejLPQoKep3J19NUR8zM6VyatLOfcrzqExpwwIC4JgjraVc70IAgMWv0R30a
s3gZ/vUJJKJKUgfbvtJWDQJZ+uUwdQaIB/Z2R6mvPJptu/dnQt4xVeGJUwEXS0J4
7FuNLfkHh6eQn1HFGqVMOuKUyZXdqPAsALxBGiqQse53sK72PYaFWOu8OyNqcPxp
9O3qXqZ/OO7ZcY0Rmyx4uIcXNRdl02vNfngLd2BRBi4UfbsLSAXTlRmM9W5qYNRd
VeofmwGL7+9BZUQYcw2HdCg+RtUgIND/X2yHIS3LENEP10rB24qtjWJmE6W45lTv
IdTuqllTr4QvdPzN2mG72tQU5cYSmYVrOSUwM9sa7sNE8uqaodoYGD5yqRIHkG4c
59pP2CXrGFdup2Zbl3sBnLU0ex4vmvWjcU19zeAjsg+rLPVHTqte68sWDd7LE6yG
SJAJdVfUMq7clqlBAqYzm5kb71uTc2O9GrBZjDmiufktWM++pvWWY1ms6Y/2yPBv
5+bdW9BgyEbUWVj1QKUTCqp/oHEWhKmW7BcOJaZTbVH0OXSzMx/ZEIfS34MOlBTN
lRUzNH9JGvdHsa3FEPJdAlRGpw0VzfWhLmXf62R+C9JV1fJVJKajZwqpYj1PY5hO
Jk/V96460Bgf5rb8ub6sikYhisbpU2BW6qBVm1HhgKzmheW2L55xTQ1LppoXWI0z
/TmgGIx1vnpGZKoi8YbHh8605ASXxVp43B11PRDU/if6VrFg7yZHiGESA4OMnSMl
6yvScQ51BDadNzUJfldPSLswa3MtM2S4EA4VQBoBXnip7m7OIW2IElB9nYNM9Z9t
bwo2pGBmK+atW1RJ1QA4j6kPjJR326JxWoPRUkRT9exM69TfIGXmCWuoPye2ThYi
MDiR1GcFPXmjtaICe9JMZ0eHFlh3ubirzF1T3MMXIcls0cM8WWcfh1N8EuuvBqCP
Dj6IyTgdtG94pclCfO5QUc4/ItoZCuxR5/7bejNyTUidH5MrJUbUL/yiddvyRFbi
IAw7YZZO/MbWfpExT/Dffz+uu9nxs+clGHFz1ztSglfMB5+y5aXE7l/Yo/DU7FBt
ynQrIGcxIpj7tA/mxj006T5QfWGECVhZR/tCP8S1EsHj4BxucbJ5bZopVxYeBgCL
ykZIsRVmbvHp3Jj6vWS8Lj3FN9WCOk3ee/e3xMKKZO28pki7JLULvN35ukIvOU/Q
qdwGMrBCgcjx5CM7Binn5CFwU637k71vJdxHFRE9uknpTeVyXL9LFNbGAtGEG34P
nw7sM5Hl8YvaUm4NLffiFhzkvwQ5gYDFsdYgeAi0h5zzPjJvlxZw+M3gZaJIauxL
7MAT9w/LBoou2HYVbOybWtS2rN8tL2IGgwjscSTv3wDaphibKK2k78JFRdF50GQM
gIWFHmBMV3DFDc+sBrkCexWkLdUxlQrUQh2AAd0pjAB1bsCEF9z7kW5AOqbFnO/e
M3o5r9fDFcaryWmqS6LcJ1o95X96z9Pk13p+GhTojZdeXsopDxReKTa4l0hkp6Qb
ZoYRgNsbW7OIIakUNgD/wHdWUTJBlpWdCirPhrLGIegDPCBGofqJkKNYJrz9f38H
nrbt0eik7LI8nWXbKjo9h+0SzfufLttnaRIR0+8zBaJyNF+X+FDDi4ca7CKah94D
YAHdykWBxxcAnCNB9YGNbIEgxI1AZnAi/TpvC8P85gKjcOWYVEzPlZhxnLvO5kze
HIEthMWYVjrJTjf1jGvjjD6vZeiksdkXJqeO5VbGnpR9J/Jfsk5x2jA2NNpPw1VK
/kwLUpeD5qkNVaZqc7BQKmV82TI61gA09tn720NJcMzygwtELx64QP5xCBnm3IY7
GZQ4Wkmrt3B4nxuUu3fOV8QI/1qURP6/+f7lETfOIAcg9DzlEDYAnP6qMq8/9GQO
irxpK+fDrWb1amkIBnZtd6QKTqC8c1v8NJN4WNEu2DEG+QFR61Kr9Nwmm4QQTSYp
Dn2YT73/vM7/nONbGY8qw9i7Kukd3PF+/BVw+IGi+MRrjjGZQ4ZN7naTohGaduRh
CknYBx3bjHKncAP85UylvCH5ehW3EUXNZg39jLIb9H0KdEH+EpY5NL90Nr4fJHgO
4dVtHcMoWv0gikf+ibOHQblTq8F+ve5nGTfCOi7DDifvkR4LzZV6EZNlhN7if2eQ
OdKIolEu3rNyoiqopvad372GIDLjAGEec3JpJ4HwJoRTnCqo4TjQQW99tKG+JPEF
if5iIg6fERcdiPY5jZGeABGBK65smHP2vCqfGdcJE1kewiAh41AqIZ1xm+SFkl7M
SjhJSLjw256LYL6sAqGSC1tgcJkj7Zu7oX/59q0adEUVqWFh6JtRk75tHpU8VDM5
mAsBrfo+naPzWD2tmpn9FzNAYodNGMHq/eiwRSdsq155oYeE6M31h7gC6f/RxQFg
cI0P5IzzuBi0enkcqcp57JGT/tWQ/iXylWdKc79hqRi5j85MjA4bcd0mBamEB1D/
VBeLylr4SeFGefMHsPpGGxz8mBmQc96lB9NIhRIQcwCcxqQ8MQQCkc4TASbzxihS
MYXf3jqsuMMXvwpkQ6JkSk6Q0ytnj5+p3nlno6KipaNMPxdTca/9wJ0eaGuQ2j7b
V4x/VahkrB+BD19CPSco8X7A8bFyVWjwXIZTVeJnWNHAQVImw20PkXCXAOuY1ADU
mtt5RcKH/abxkF27UobY7wK+aDQV8nIvmIxfwBrkmbqmkXmaFCiQHZiLyfFOKRvl
LVPHoDql9gGWOUsn7hOIZWVWuRF4t5AvIE1383O+L8retbFGHtX6bZHE/nC2gnT3
O/ohsaXHSMnC5T/uJIKNH7j72XDoTm83/XacekkNRNpDcpdi8mJcaODvsjJSvQDs
OZ94vJQYvkZ2vQOo3RBAcHqSfidvY2wT7Z0MJg97KrwOjr1wmxxxlErwBcn1BkKT
TJvlmeiTUR9S/KPf8kM8WeUJG+rRo6D+UKTTWtGZoTdkIxzuET8go9Q/5ekeIOWw
tVrjM4dMUPZmZbZACWUHoIf62VExaBghg5Eg9tCIW56XzGxA81iyBBoeIlf4ZVSG
abq7xdJ94pFv2GiyIRamy94+y6RDdSpPH3ukKsP8QPsL2Q4xjHmA7f/Ivuq3qui9
Wp0eztuiD5YOMFReNKm5+wjH6sRrZlPRTwbbdB/5jAcKsm9g+evhgfmipAwDhF9H
i3OfCfj0ENN7l5xfG3IQn3GfrkLp6kifzNHAjn28ctfmJlfEvF22A8TOHF/FsLk1
9BsM4kxZPzv5yVuB8c+e9lCzltg2D3ZVTrdd/x2S8/EC86Om37KJea1BCOySFcUR
pWWpv5GUHSlXkJz1k6N+71iwXToIrLH0Th+DpV5Neh8Gbp6NBTsxiOGAUCH5dHyF
8rkOFz7fFsiKbUjP4V+yGy/rkUf84EA6AXwgMfS575wFtKTAffO2emCYPIvcC2nc
v/QpZfn6s3qOyAynjCHd94L6TuYTtRdfV+yzBu+cP9vnWl+CCYQ+Tf9pzLz42n43
Owa8cKxXwkiOu7oIxjt54IzcogU6DEUfa42NZkTuttadj0OutYa9rFaSJtyAz405
m8XCTNJUVmJntDQUqchyq1fcI4Mzzq4P5zSqskfrO9vODOHxaLMgXvZEiNadb855
himV4JHYunFEeglTyPP4jYifCHcJzRXwVBU+d24aHb5CGHO1ppLYYm3w5gqLnRDq
OSmXInLVES+1wpQRv9A349gJ5r+ySDiT7LYI29Knd4vPsqX3gMM6ud1V0FfWI5y5
83M1Ol+N+Mcw5YWx/rRCY+1iKoFXRJ+J6JRsOGUAs+EDhunlpuPqoo+BLtX6XP3t
mzYQoixE9Y8MxrpFQuwFM3FcODfPcSKk+UN5EyqXXbvlNag2NUxvgC4/kgRXTdAP
VxlzP7KHIYpyqUTEzn7ZSEuwv6fUc9mFKqN1hzoDxsXSkKw1amFsB/79CULKfDcK
ktqslinSwch3e2NVj3Vb6OViP0mioSD1i+DDtdmlprDCybgVAsj9WX2E81m9k/9+
CyPkjPJEUi8SPK7hxHXQQFIewiShcTEhaRglgkdXaHYF3ctNiduXmZjs8G2AfHt9
FVUmdroITWvsnEIhErg4EfqOTvjcRzp/bOesC/pgXeK5UfVf6NFlX+cY8yEVXA82
CN17xw+Fr104we0bfqIproMOxqx1dQnBRvZfZOutXxvqblE1kxdKOVxfG9A8QKYS
PYsxtnZUXhD8U/97neE92REjz22frR/RdThJpfk/FjTL1AaQo0T1xTa3WtWLyuZv
e0YCTezxphYqHnysuLKKQaq+3W5OnaHRJYVepgfLWHkplSpabq2bt8n318mpeOtB
S21jqv+KBH6Ez5LtWzRTCuUUsa6NtYwnk7C0MtEt+BU6x1jJhHP3BGO+ss4xX7JC
kq0pR8QE09bsTvtqXwe7DyDwSmduxwn/SUS1CCevHliVuXuipfXkbSq/SoV/A44J
9SXHEacDt9CH7ERRFlHiTT/D9jR2CZ8rESbC0aHkUnFsizswcmppDxyQ90BFKFb0
mRwp9N1ygF1bJEfrqEnrPALwjoN24p9uRtPWsiDmZ6myZUFFIz73R1kj/xI9zgeN
ml/WUsBEpyjsjT10VMPKFWx+TxOkyLB/r+8C1nFiBfyVar9JkZsR/cCM1BfarM3s
HIpHhAH8xe7+r7brnadJIx/1kjuH0/XMgE1fxvyKCrIs5Sc2pYlNUgV2k9g6L4Hm
fVXoPX1/JW8K4iFul0riqReqPMj75+dsS0oqu3N4svnHEA0LUjrH/GtwH372sHB6
HdqS3LcC6+SJqtCmpmDbLirNyp0n7yHNy6ofXvEGhO5i8EfTiTUeI/XReEQYuKVk
h9Q8gW4YTaGYXM742csZRYLCXhfWNrOiWhZRM/Z1D4DWyWRIWdGFf5fsBcXTvHMn
tzIAQqMHabTEkq6v8m8IaDsrOzKIKaH06pTcWo3OYzy0OqSr/Oyqs09u+m8rFoBF
C9zsJTAUTHn6Xfj4dUI5LKPJfGO5cVnlDB7eYJfx4KC6mZl91daRdaCi9jGLqXgR
2V2cErK8kL0b/i0CfjZSo3PTdsbbpbCEa+3rTwdOyhPria/YiOHdwQrZOSVzV0cT
CgHABA7jfHnPy1U5zQSnFgEkpXiXoxQ7c9x1ESxnxsXCnP1STgIyDE0obpsj8ZI4
i6jd96cY8gdut7YHt3VbeDOu9+fuTw/lwhJhYx7JbMUpdUcrKN/QVuJ3qPV+8zZO
dooylzkzyhyBTY3opkTjvQOdj3/tBY62vnLqdpu0otgvOapN3g45ctUxsCqfndBn
m/skCuF5pZ6P4VhQ92yYZdo7hnUU1Won6dQZRhQBGiK4YaJYyUOfAKAl1bHpe1Xx
XScoMVnP1CMNlrntizJ7QWjawH5Rxb3NoxdULyTCpCfMcBQ6f4jxCPctCBGQZ39d
9kyNu8mmAm8xrr5bcp45hjuhO/ip0HsFTzPRqhZJeA0LbCxPHt7zUdJrMvFagypl
jGQocmu/ENi57QPGGNHuK0O9bl5LBVMatW36HWxIPPVHNzkTW1wMsfBiWjo+rXXm
Z6d1vFXC/gxuMeTWQN/lvW/mzNLvHkx/jj6M6pz+1oFMZUAU0LP00xbbX529r0q7
FTcbPyybIxjZdRfQIWFJV/wxt8x0Uom4ts/2PpXeF4ActF6QAt0RcctldSxsrPYB
KrV+EFJmrJ0JF/AzrWLfxYXCeG1UhXCjU8Wk6s0X2xaDhlNZKmhXU+/QJRsCuc/L
uNFa8eZ5uw+hnblORJpLu4zwYO58jnJvwIt4aPpljm4iws7fD83bhTI/Rj+/Eyfu
4AJu3IVZ/qNbxHXTKjZqNETMWhVix99y0Kg4L9qnWvaYFPzShwZVkuXUhv9bmZu+
e3LuLzw5wlxYW5l321xGC4Ppr3re3jiThWUv0C7cAftqLKjUJE+eGG0LvTEKiRHc
XbpSZGfobuJxQrSugy67X5sQ2/+CMWWxQHtPaQHljDOGnVks/4ZOq5PDu9hHCBAT
OE88tm5/TikppYi0Fyy0kepwnF/v0PbEa5jha1aR6ITZkjkxXdde1VCjWZYWr9Lf
F1YcGV3v1JVUS1iROq3NfrcQ2mVzbhHw3AxxD+6VdKaffxGD9YYXR/X/e2P9kYSp
uita4IQSPXN574XlssnmZ7gftMJkJb3ig1piq7Gi6qBQKIorQGe5a5HAIzJVgfC+
WVyeNi3dqvPZH0rXU3qAFNKGRFlwaHT280e81lphpXMgRwX5SKSHURjQFgmgjHWt
+OxS/LPcawW5VD3Aj7wvt6+Ka/u4Wntzl6nybd3Xp/bLggPvBsCDYqr4DwS0I1Bd
tKholEJipTOgFmtn2hVrwDYjWLfapE+CR0iR55aRUx1naYAZUmPu2J2p87ZHrK3k
u85x2DgeDKOh5/cbKQPEXugWeqenMnYEU53GZo/4eE1IY6mrAi9N+TEnXJ1aTLKE
a54Ym1gHuv69vNCpzyaoSgU4Hxb+f31ilTjotnEaPGgqGMFGLpF3yf5mWzh6uYCA
eF9jRUngkpOuNibvRLW1x0CTp2YSPpJnez6AipFORAEdkfuA/gTT2ABNBB7RWpIL
qe96Q6OX83jWvrPiJBTkM+JTp5mDA/KS016eFQg/bTI8d/nnsSBAbY/jyrtol30O
LBVoUaB1ynSlc01OSfNc4USO9Z6Z1nYgQTd83uHw9E8Azh12WLUvEfpIfyMOq6j+
+u/1wZBI/kcF2fw77VzaEO84na8qMzNlamX4L+jsOM3ePlDj+fp1NvUwTtNYHE0A
uE8GIl6v7a/W45IWgqb5IhXlj77jax5jPMbyW00wY1yAUMRh7SaN6VS/Y7MC5vkY
408AxUdoExjBO0QoFqiuG/UzZ45E5Vi3nWoXsMwrP3TlrQIBxbpIg5FtgTF3kGIf
yF/+L75JQYMcjWFuV629kA9jwZVDt9EpAAP00nVWTSJCcBXRdK86kk6btMq/Yjey
FGJXxhieE+qEVy0/tRoT+h5MkK3CIvjGDGIeBVNCqAfS5IYcVj6GFR8YJeUN9Xa8
0WlKHYY9xATZzjfb762ZLIwsKzgGaVAOU1my7rqMXloXxV59dI47HJAsjCO2L2qh
MVfdiUV9h8Lee2xYAsq/Vw==
`protect END_PROTECTED
