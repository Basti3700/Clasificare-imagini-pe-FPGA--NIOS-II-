`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkH9Z7Bd82O6425hoXDMytv306Q3vp5p2JI+KylV/7A8ZGWnbIkRc+PfS/G/wDbj
bRclLKgLPGOJAvMx4Gjfzwq382TQ9MZUofD2w0HNnpfhLIvnNbp1taRtvazlNzC4
4uDaCW8xwM6OuME5cRNV7hTgoP9fV8SQDfy27Hi3viD0kPFEhSJBCUqEitT/axo3
iGmPPv95cGudLMzKAp9cJVCeDEjFqlfsH1OX/SybepAYWVUTz580GvnopoJnQhrN
2NS50FVl3QIOOqUcHwId0O2jxzGjIWJZKbK694ZeHCm0NrbcHhAWjXVjm70yV2at
wZOXAtB2DS0Ul30sDbIeS4fuaxpmwSeZJN0fjMCk3P2VDdM0POvC+OIEdjHsICcz
9QMItJPz+RUpZC5sr469u4+s3EYwjwrFFRb4GiOcbYAzVh6eMW3OdwrxdLzXLTin
rxPAQc0UAGS0yBLeYR8hsfDu9RQkEBeyo/512ZDoFupsiI/Zb08len5YeyT07Ztt
AFvAVgpbuKU44Qshg9fERwL9rx51dZ1G78LAES+pOg0ZdrfgeZYPyXa+dlSzOFSH
tIDtHHzowlCBMuzJLrHjNnGD1j9GGtPKlLBYq+Za0pwVruyRRAMT9DfZxSINksNk
WQuU+kXiU3/eyRa29sDE2sDPBFG1Z2yjWxMeE2TSYCrJah4YB+EZ5SP8N/D4Z32L
5rwPzwCX/5Cnc1ibiaxrmon21H8A4F50Amghbvb3hQI/KWE3A3BP7VdDtP93c+2+
3u+Ibpx43WbiqZFOA5iQ3wKaIv/+ogcy+X69Dt3UzOBqTGifcutYUaGlYgSsVXhe
9CTS2rTU5vQqh3ce6FExmwQH+nN7CLrCfFC+B7FXAV9/ZrzLTaxptgx5f06bOknj
Zi3VX+T7aU26O8nN5z0DzNkRKSRo3UDA4RE6i5Fx70nJhKPtpa7cKjEAsZZdJ3Z+
SxleBDXlRv52ga+AdhnQkNUJT59fWugeWiC3DZZglyZRAQvy/Jts3RdkuUJY67ig
zmbTA4Qz3++yhmjfbOM+1nRYqeaJRyt2JoAMaZOJEeCC82+kn3u4SKIaorkRBmU+
uVYibkzBGCD/d2X9W6n7WWqcmqcudknhhhsbyQtIthfr+U+hWN+roE53icNUe7BD
D8SYPwFtqyaGDgD8SDfLRIcmI167dM1VHZn4HGR1BVxIkYsh1ma7UCzO9zyIQuZt
ME24gLl814+JAru+uV4WAtMcw9+nFHyu4NLnEopS2ya3L9bW8CvVpgsMGf0oB8Q+
IGRRKEoxop/sqwk6L1CKPipKNO0n4LQC4/B/JpKQ3bfLRq/R9C+/QgQhRPEeM7YP
BIC/Lu54xJ9Q98tZfMrTK5N1FqsadRpkM9rV/bJtPXubldlexmOVYpUnNPIXLfzA
z2fUe55J0I2t9k0WRqo+DScCft3xfcr1Gr5eB0QdnXwn1mjJxB/LyL4tbbcJ998b
WAoFmUM7uMy0XsyIUWCJ8RtcXsEBK1zPTizo/tx7v8J69xxFNTVDBFEnbu2QK3f6
FyYn1wWCVFtfMNatgOWfb/AdvNNKN7ebxdO569o5gW5agKtLeEddMja/g/wll7/y
rUDn0cXTMYz7SpOfBLlm/53LvNWHrvpV+EFz731eiYOeBfiLctLnWkxzEyha8nH5
FOtDoN+JFeyapMudPkuPgayyKpswnMqkoQEKmjifvu7g3SdFEDm9LtPvJ16GcFNX
nHWzh6gUH4slKB8Yw6pbZkW+bQu/xIYFUI8vy/OiIFDpJxk6op3d28rC+Y8xsxgn
VFe9A3JeUuu7XkLJndtDjYUk9+gtbMH8pUlivYt0iEc1HUlGhCVlboHWv1bc1hO1
gNZD7r+30YSZgXFPpyb2u7tZSkmuocTBoQrVNRbHDpmV9dqow8ecTDFXThxTluvK
lrn62s5cv2WJ30zmGEeXoiZ2pbY3n5qVMSS28H1e9SYZTQ6IRoiuKIKAozOTiTC3
UTpYTBosrYCY5TiHIulYTA9YNFA9Hg0HCgM/tpyhXixMEMEZTG0a1dLPzasLgFwU
eYFaJDfuHWBFpRSdr6zjRUOaroM35+UExpM8dd+/3Rdq9JnxO6hED+r0Jxif6n5j
SL3jNkWodDKeLzjo1i77wPNC5uGsbVrwkjZ7D+a9MI9IUIAZnkFxRwqoFa5yt3cG
lTvmtBHPYk6x7rPbXY25RBWBK9McgCl+LaGgONgrM9onGDVkQIKOVnF93i0W+/OL
9JT/lJgSQX4fGmxo9zWO1tagZiCboJu3iQd8dtDM2Xor4PB0dx6y8HFjBuLnyr4y
ARFvQ1l1QGuV+A5EcxAHXFP3gyhUcrzbfqjprEOFPaGgmJn+kvnm/wVu66QIVX9s
mELgS++r4kKVnJCbyWpeANmCD6U4AhGSUHSwS4uDMCrQWMudXRq4g3xWw/697Sby
8FRtZSNkl5u17+NKm+PGfv65UHUEQ6KADB/VOnMp0qtja//z/9EiXcF0YtLhmCvc
P8N/aiYv+r6HAz9HB9obDJb0BmL4Ucr9slZBAHj10KjVCDgVi3p79VRmJFtPBevz
veXqV+7dvOP56QCUV5t2++Jkvxs2Nwum3MxswgwJV4xWDvRMl+eQuRs3kkWJRncL
eRQNLcQmYCVYA0ZwJzCcI3UQ5ZQRyTWQdE3m20KGxdW8wrjfVTz8jRNx2zomzqb0
C68OoEdlJ3PYUM1BX8qmnxVnUG7o9/I+yqerQ+j0oU1yiusvm+fqB7/O3xAFhPtW
rscShuC4gvCNJO2ijk01QF5GMC2tYzV5onfssqRxwOrecz9baWSFS3bsAhn1/fur
r1549De41A3xzLrJ9C32sNOX2Wu1055FXZODElcR/DxuzDAADkOr+9abe2dQMVms
J4YCyan0FqA5TwyuxHotioUmpHnC21rjroNxccPVFwCeZQH73m6zUdb470xaMQxY
WT1REr7KKhwT0oXvJKYUpJMRMLiQXAX8x8S9XUzQict6L7eDwa3tjQHUgFsb+8+s
fali5M2z7lKUaPCcSrocwDwPM4Xa+I5c+v+GZs5/PKUXSYNLJrBu50lVC/cNyGNn
fGWYJluhAGs+gNjdS90ZmTTQcFhGlBF7GsJkKjl4t6R8zTk3GHY6+DcRNl7NOlkC
50nkF2QLC0fEjEhx82+faMmgERxHPaMS0Je4ipWzi0GHpRtf4lADGefTSpyfyc01
gfcJ1pMoDPdZQYIHnTn4U7dViaAHX6fiHOhMZV8egHi3VrzcP2p4iNT9XrPnzgrQ
3/p/zoZdO1Pkg49zq6DM92lyEs6JzDJFyVqwcevk5zc0fdUvCUgNZCbmqWoAE4ir
WfkMpOBsNFJd8SxUXfIMZLt+51Z+Iv47NqgO6E5cohJEwsNaVECNLEzfOusymgi8
8HJeIAzAfXG7SQKR/Eki62aIMbIK0C5KEDzJraUIF1YkL7oNfVtqnsoY2aM98q7D
x7jWD8u12SIfEEgddi88BqFaX1g9lKy1rHGDlaZRpjTnK1v7NtliMnBMabC8m8dL
4b1ehAo2CD4nNb+RKNxBMTF7E3Xvhc7WFJTtzGaAINhyXBYCmY/+nbCBGovG0FOP
DjXdbuln20hKIUSS4Vj6cGweUEa9JfNk3ZgE732dIsTvm4eassRwW0YNQmGyGNFY
Q5ZPvv1Ir94Rbf7dVipvg0eK03IvBUf3dFPg6QfqMkgh7V4Ks3vAdgMXaBi5pV7Y
vx8e5fgXVIKFBlUEcFFb9Rqwdbn7wHx2jMem/kL+8j5GzvgYEcRtUhYMTw9WUDOD
FvwBLgvTgN2vGcHYPNTw5k+UoPZ7pm1xKHPJuCPHPSpMU413CWSmQpz7301N3gfc
nTGzVW/MqJUcp2Juo0+HNWdac+KoLa3Mjio9XGbf4bjKIHOghw9qW2tIlIe6Utl7
Gcjsb866QLi9WIMWyph6P2R8KJmML+xUlrVOEbaRi/TZLPju2Fu81DlBJzgJCgWn
vpjR9Blzgs13/sqCZzoU4x6vtMVzJZKTzv3dbf+5AiOJ48SW0MQnM8BGdfDh+Rs5
CXurzW4bDOdT97Iok377MVMGK8AzDIVREUHpeLrttxegubfyniaUMnOg9J/TQR8E
UgDvLJ4g4J5xZ30Hv1haHoKCz2VcNruljIUnScChx8G8Y9F90K8m5dHBj7SFET+/
AkH8LHS/XnAoHXpN0Jx1K5yZ/hEpQ53CQQSBq0oQh3sQ5TaXdHBP59PPDAsiKGou
HhgMUfnKMjgYwMsdKC0u+5e93b+gj/jGk4wbQlGlfonwx/JOobRKuAXUcl/Vi/nS
hol51LrZ81yRbzclyQ0SqtTIYpOQM1cedBxKuvHkvy6yAuv0JkC5WL/bo9qEvJVC
X0cH09pSCkaHeUA80aMkvhwzmPilGaLGYopNV5P3EAz9qAc1LJkygrODR41Xb0DQ
`protect END_PROTECTED
