
module ipselector (
	button_rnd_export,
	clk_clk,
	seg7_out_export);	

	input		button_rnd_export;
	input		clk_clk;
	output	[7:0]	seg7_out_export;
endmodule
