`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q7K1V444rNZPa8LM/ZGKL0XeiK5VwrGfZvd3K/0HEL2vj9Rggp2NjZ8nrYLgOdct
J9DquivfIXpfgmJU1lxclNOWId2XDAXbqHj8XP+Unb2FvQ9HRWWV8IczhC3acdP+
lYc/wzyT0TuOVV2OS00oeHmsG1uELKwEQCuAx6K65spAoAbNFm127v51sBOhWz+q
AQOMugJ+IekjTOZazs/5lOMQZQzSA0z0KJK5yV06WpAv+g42RwJfi3DNxqo8Awwq
`protect END_PROTECTED
