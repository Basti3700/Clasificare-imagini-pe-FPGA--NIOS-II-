`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GFgQBVo89CNM3/TB/ePbaVb8OiqGeYTrOqbmaOErFMrPpdUnYawojbJahBAUGxg
E06ou59fvVDqePaaNLpkznulEDRfmH3TMlAU7+sj6hSLC8xSsagbC9GA5mQR5mw+
r3BPkv7AUDGJCTW2zXhcJDO8uw8LJniTz33VOGiWvnpravJPvCithKFaCxbxiYIT
eaHc3zpPGF9edeUNQOMMdpAVQNFhDcGYEQTBLxqGz3LLrxnqcmJtyd6daVrT3OEY
++OgSccc0mnfzRq3MKszE0HpMnV10xOkECHmnN6kGMHCuB3k/D3dFAz0eBF4EYt/
67NtZR3+zGLZr47K9TH8yYYANce15U1snTtxd/YpwWeFh3l43Hh+OrwMlteiPrLS
PLqjAcCJx7EHW5xooh1KOW5htdS7tOSgYtjkJZekwGJJ7SrU+umq9Dho2+r1R4X4
QdnbwM7X6VYn27EF9q7HVREuoakqfUpRKhaP7MMi5RgO7GbFrrJsFgkOgb6G25WU
z77PTcf5kAxWO77g+ECZJma4oJwnq15oY75NFHyTYUIG5X5T0b2PNMV8S2y0HomM
g4ZiO8hR691eNPVAdIL2LOcbgzzRYBd4DxVCkM8SJwDFaOdD1PM0/EzP9QOyw8s8
cgNHn4CieX78YXbwBBN6wEILPL4qFQr09lRVm+A0WNV8J/VRTRZj6Uoxd7IX9URy
MXT29fVdzX20tLVw3NRxI7Bsw7ZyorxpZJ4kDgvWymRk7+Rp2CjipkvxmCAdq1e5
wxv3dUFMvjIqePEozUCdtQY4smhZdul9an9ND9bTb0om7agA7YsJG97ygXwaopBS
`protect END_PROTECTED
