`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FB1fJbQsLC+00nfrPxki4jBsne3kArys5ZoaCt/OxE4XRiRf4C3k6eMMsYL5jBbY
cZHueo2xaV+rKL7B59t6eSOuKoSRsiuHjmxlMvNk8Qnm/fH350WRg/QC3RC0dfde
SUUOhchD9ZKhVUosN7QWqHwmIKy21rgRJUIFNoL94Pu1E7np87P5pkB0DTXCpVpQ
vSd44FPr2Z8CHkCxyl5/E6YkU2B8uOoJD0uQ3zx6lLdJTUGNfaGsTSgOK2XDryZx
tdBKpbSU6TXrngyXWkfLj6l/xEnVCNYTN3mRll0RCk6Wy0TWBkxX9ud9aTuHMy02
evAiyxrkNbNXLuUySWSBLAJo5Kx9Or7ZdFPusP1WwKDrmZ6SwjZXSZZxG22DjOIl
qfcvZGldy4eGAulqipT5NeYKtWB0mUthy56AN1/ugsGX0leLPR05/Nry2a98BCJG
7mlMXUV6rrQMIdWn3mGRgNWhQKjbznKBdMxvbKY0jmpF9Ip9UL7BNnmewscfUTXq
Mu/eWpR8vBdk81alpDGKCcQJi62RYKswN1+kfQ5LCo/RAlrDWQ6u3doCjFFEY4mU
onLPpK45YYFm/8H2do4gtG7zSCBnUpWV4cTymBPD4YUDQMl9cNYwWEAHmEweHU/7
zeE8lbOnHKJ+flbzJHQjYf9f3bv44W36PkZju/hryirSkH82UE7+STV5jL6IB7WG
MwukhwDC/jb8hT+f5yQ5Zy0T3CE4nq4YXn0pTjK25hHBK8sr45vFhj6ZJHJsXpsH
IY8HJ4SJT8i/3Kp5Vvh6So6igcctVveljhCW829n5853gTQEUWGPNYSD/g204Bep
ZGDW0Mg7pBrxqaP9ogcZLJ+AJZX1B++hQNYPqOCVU0imgZquL8afebmJr2+dDRl1
oTnjgvDruodRwLsKEu9YmBWn5IA39YXL/J1LgsSpq8njUqC5OwfWIYIlUvYCOjFY
Ve/T9m25Ehex1eNU7bteY8/xRo0V2RRQ+7cusQzWkfU=
`protect END_PROTECTED
