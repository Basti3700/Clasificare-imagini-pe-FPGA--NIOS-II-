library verilog;
use verilog.vl_types.all;
entity TOP is
end TOP;
