`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rko/dohpgXuKmcuXgpREOWBTndNFAlSzbkry8xzE+zlewlEOHdw+9KJi9Wt3BxSI
yCIJT57eEKYmQPyWc3gbRmK+A+u9DKxCiXm9uYausNUIzfGKHrXu3QmBsCvjjWtp
KvPnWrmks6Bqo/5iC3YiDMJmdxaduCTIdWioyVNrz0Od71A1HfeN80R41qIhFfVR
yAXY1ew1PG77jfKIMJt8dAHWcLup/J7llZVk0fr3TJNI0hTSAYp0BYSG0NWKcoug
XLTlt0holCD0MCgWn2w0PPDnewbv+OlbRf1jzEhAOtOFGDsOsqK/hsh297P1pkOx
R0j4IYyIGt3ZhDLwRsTPZ4GytGXfKizNncrI0RB0uwD5c39vAcL/E0YgP7xaX14d
w+Nv03eYQcRJEpBqEa4KRckoe+ery3bfSIJ0VZtZiRFYVixlbfcdc0EcxOAxHl63
RDTH3MakFBbGoN2eTJWKLbzsjYA6LRSlo715thOhUoOyhFh2LOsnXKcju5/f3y3D
f9kjCL5QeAjNBW+N/qDPosYrLJrT9FcIomWmLbADB7+NLs+cHyAV1woWeCefiAcy
c8RnJGdnpsquA51K7OTyFFKo77puQtVawuYbjLjrNlYGxqFfLvb/5vVPg9eIfJKG
tlhdalewhVnyqL5Ri1I89u34plBm4+s5R5zUQdkWkPOh2vynpkm+xni9aol2KSKN
5iVB5kkOFPe88UtChi0IcaopdCAFkV/C3mYPJNJBVWoRi+XrUnmpOLTEsxaqco3Z
E8GrbUFBgXwlrLHh3/pyDeSa097SJNo+p0rbKfGHetDD1il6qtItQIcsJAiIqIBk
YtEQFW3gwEHj0l/MfAt5trMlCBaK6o+kPojlmXqI2XysT4k1SMs6FsUhGvAeFJ8T
kFW5K744SciZzz/VqJDOI3j47bq7E5fJmGu6YjLOQAb4GekYOIp81iMKClsYD15Z
SHNx/lpCVhcM3pbF3r5OZEcFZWxjhwdkJbnm3tZsQ2DcTcAIq5fX/V3eLtOoe98t
ocXlTitsIBSj6A7XCVzOUnz+lu6tt1XYoQVB/jHMDLa7EQhiIas9B1ZaWgXCXIFD
h1XtGQMudrp7x0RHMrB+IDqLpwQ9PgAPNQuJ4tYGpbwczrnqDBJBYkK4oMRKZGZw
7IUB0lnJwP+zbW4aVG19UpEkNdttFrDkGX0P58zRMA39oEoSubGcyVTb3G6FfQ8g
CkXjFs/8lOdzdWx+a72k/Af4Fm7AziqEYzZfLZwVR/LM5e6HMHWSadj6XzWVvk65
CAEnNyUG0bt5HBQnO1MYTg62pi3naK9CIP++NB2UVhs1NvItQOk20+ulFguMGVOu
o2MaIp7FViY8TZqikZODr7060nKvI0wJbWlNgYeBtkq+xSHxb7qpJ63eWkj+eFCc
NcaxtpJTQU/eNhH00EqcYxZ+LjSK7MdvNerxr3cr3yGAzxCs5Wc/fn6a2LkWXyjC
yO+vO+s5IVsUj31VacfwVHwLcJwyHqCy5qNw2jDLkrcXq+fPCuIq+Euw5H/3shz2
eUwSQ1RkXs8p1gOIRMIMNNAUv3yfZOXa3tYhp78Rp1CDhe9vVOep8qNyaIbKy0V7
xA+SGKvjcHnx9y8bPYKUWIiLmZ7CIXAAtEtulFPPuLD15F2+B8VC4+ixyhTAIIn5
oSbRDjsUSSZ3mdMgSW8wYPVaeIiP2yIlpdzb+YLTzlCrcOen/rZ1nmzdnQpRaDtg
V37AQmCHDOcnel++K642BdzjMG2CtJsg0cCZF9Ek9XNw1aYbt7TowdunBtw/zBxS
IgB0VOAcutpp4iguDxjo5+Y+Xv/D/Y7oesgAQi0wAeI21gXXe+6wfTuFZFdn3GmD
HGexCT13ryR7EEr9zpZ1MTeXv3SMdQM4IpI3NSb+GlrCEbLHmPJ7bojac1xHlkEm
wxQtFbSBHfPi6hce+YqIPVaE8cC5EDjWIg9knvRoZZOXQVN2IzwwzBI229KzBnUs
g6bVbbKNw8pZWbDWemM1POsmJmcxJU+WZO+TPknQnnF8dXWUC5/rWsMZPx44rF49
AocDmEmr5ZoLcqJF5ky3yF6JKaKqfINiemz6gTIq2YN6wE2rrGr3JNDFVDF+hCCS
sE6wkhorUZwAyJgNqJdjOxA6H1TsuWCUApcGzZ0OQYLzYPbTyG5+kjN27hlkcb4p
F6dweFNPI416jbOKa8lNyKTB17TtHpsK9tKKEeEDukTeSvXIwtcn20WIv0vb9hn8
muS2bnQdBcn9NigC993IZVvF6YtIg8Fdkw48951SiqfqSj5MWDA5nQT21dxkRJc1
90mvCvgI6B0VxOBTby7hFhGqRCSP0/BERCXxPeXUV+Zl/VEc2SoJ7Q+F60FqHhar
QuEip9XeSis64NmY/XxebCuWjFUffbbFLiRpPL/3Dz8lI/Vepg+rTPfRGeW/tITo
WSzv1JqnIh0fZdg51DpyDgv+k0vhk4t9v/tCeCrW0/dDf54ZbN5F/RwDQ5dyaS7K
BDZ38lMeMuWjAK/YRJMEKqUyuP5E58G+MS7TRLmMkbZA80/oI4JZ2iv4WEI2RghV
HtpIFy9tZhVVcrer2LIqEWyaO3ehkWYk3f8tkbdoNJfgDiB4tSV/4j17R3intRUq
s0l45vyMYZ7a4t45FAdDVgMjCCkZWe3EAwTp6v25zu3YHdq1+ToQ/kSklQg37K/y
hpkBE+h7iGbUOq7ptF+9ODpqPYdcXtb68G2ckg55zSQm6jbD+P6hmTWwJmXJO2wa
Hin+3/va/JsUbqjABv+Okj7faVGuUR7UDOpE58SY55oG1Goo4UNnzDEmQ62SozSw
PhpO3WHBWf34wtiFfrPRoi6YrWdwXcCBxW1DYqApzNJn77Nfk/X2uVCDU2gH5qnc
/m2BXK3yoanQZW/lBX9SVgltGt4jfMlJ8cGH1qZoNMyV2VTuSOEjZ4gcQ/HPTtm8
MLZnVvj617VRo1s9RPofVGYU6D4NVCECo0vjbxRsY0uoQ0jMflrmW3/QGvS+hD4Q
jimJbHfwXk3enbV109xu52DWJ2mLpDLf17NZRDoOCazBdzMbpF6Ke4IeHLLePe/k
xJJI8Y/R/I13qRCMJcKivDD131kA8bENjWu1voeXG3Z1UxUwCCi0VoJ7qDNuAxEg
berG3jNBakm5zI8QDrTPpgRo+z7qfDOFQvkUYWks5EIJE5lL5VgZk/vxP9H9w7PJ
64GBZbAXIguYFX4lpkwfBHNNbZii8onKPP2x/hN5GXcGyRhfzVBAHmcjwTUoSxts
Oe+K5LC8hph0XxghASvqRSfIppoOCZZIUTslKZrIXJIawhF4+QZxIZDfGyMcGfy8
f3lyBc1nmz6xUiFZvxRyu9em3NuBGjn6koipbnJFHY9g4E+WN9FHsuoUuGdR7Ypn
BoBH1eHc17kkBtRyItMkoly8Xh3pzghsLo6vJtPJBErr/Lgxu/ySW/rZbnSP5FKa
dgXydC2BlK5BpgusXKEBqSOeVHVlRbpq5o0YyjikgoilUEOcx3Q3fFFRw+skuslw
BoNWVjO6STT2vyqpoH/Csumrf5HrwBo8Ng+yg1X+xLoXkRRY2VDfmfzTxFqv6a7n
7feci4xTb7FFcleVkYK/Q4aQdUR5ZNYz5jIdlIdxDAaFDcWpiyA1DR+AwKA05RBD
LNBDNYpmxpJYR44cWeTWtucXcwm5rUNruiJM8wZcPxgOoMJ7PNmlIyt2XhYp7AgJ
Vcc4qMg0QedQphJ38rJrD4PCwxN73KTUwDfoY0KIIyRgEZ2g9BWgTu65ZV0uqwp8
PnbsKb5AZ0xhpfN5WmmHyZz7D3TEqVoL/M9tIEgHBTQkya5T0tbobwJmUVVLTZyl
AxFGIKUpZi7+zJJDgP0DWfDicUbeWj737kQpDZTDMpW/PTzcSSVAyP3xFqImvHA4
lWwe9BqQGZizs/i454crbDkmssPcsyY25jcYqaK9GJN7f69/azr74dXTa043EgTI
op0L2TbEe+vRjoFS43C8BMi8le5wZJQgZ/VQ8bhMl9UkQWSiTX414ng6votulf20
0ckcvAKpcil6kvuSQGPARsI/Mz7t25N+PLEX7/BIqNqkRWgsFkAOSubxzBtIjkbm
HQbY0tAkhWizfyBUd25FbhDJ9zXCwV7+B9zA8OabUWiSWudCfBBwT7CNgohWXuh3
zJwl8gbnual/VY0ld2rUB5GewuDWM/el7M3uvFyeIXY9lZTtsiF5kzjRz+xv9pOG
ChMmC7ZNNW4o8qudVj78krfIhqH+Uw/qVrXOF7jjneWUKpuc+umY5JMVn9fQjIM2
MgC+jU7fiB6GgBGKX1+hiR2Q2OnXoxFzkInItR8gQ4SZKZ04YEI1izhhbeSXUSTa
kw5bUpaFZ5j33qUVBoxytJixnfC+lKO6FBHriz7zYXVBRjZvynl3BOQNBfJBWGu7
`protect END_PROTECTED
