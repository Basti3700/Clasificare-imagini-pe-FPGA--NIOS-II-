library verilog;
use verilog.vl_types.all;
entity conv_2 is
    generic(
        S_IDLE          : integer := 64;
        S_CHECK         : integer := 32;
        S_LOAD_WEIGHTS  : integer := 16;
        S_LOAD_BIAS     : integer := 8;
        S_LOAD_DATA     : integer := 4;
        S_CONVOLUTE     : integer := 2;
        S_STORE_RESULT  : integer := 1;
        pool1_result_base: integer := 4704;
        conv2_weights_base: integer := 156;
        conv2_bias_base : integer := 2556;
        conv2_result_base: integer := 5880
    );
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        conv_2_en       : in     vl_logic;
        bias_weights_bram_douta: in     vl_logic_vector(15 downto 0);
        result_bram_douta: in     vl_logic_vector(15 downto 0);
        bias_weights_bram_ena: out    vl_logic;
        bias_weights_bram_addra: out    vl_logic_vector(15 downto 0);
        result_bram_ena : out    vl_logic;
        result_bram_wea : out    vl_logic;
        result_bram_addra: out    vl_logic_vector(12 downto 0);
        result_bram_dina: out    vl_logic_vector(15 downto 0);
        conv_2_finish   : out    vl_logic
    );
end conv_2;
