`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Km0kUHbS7wtRlP8UEBqfSTqOsqAWHkEXbQuaow5Zxlot4CSP4Rcy54a7PlA6wq0f
3KK2xydzHlAG9JYXEiDrIxYYeoQIH1sHJBIDQjf9VRg6bHZeaf/fZH+C89VEvyXd
KoJwWO7GChsQktvdAJGuIBUuknmGZHTVQ+O62usFwTQwc5iCmqQebrjb3FZD4Bww
xvA38prHZwIrWOpgAvBFsR12zxnFXBe+E6QlSSgEAv127XwnrSI4bU8HnjoVFp1Z
+liYFDaYV24bFnvQz2YHLJ+gnVmTOHQHt07f4Tkq4oWX9Hoj6CEf6MLd4xrustmi
WSnc5ike83/HdcDn4gZeN9dQ9gAc2nky9s5QKe2MMFKucNAB5sdUiI36c73RBhxh
s4vrAV73LYQ3f1nqqtwhjd+Dqs8pBl4BGTttKa++IU7TFPyoXJhkWsBLOpNdA6Zd
DLcdb2zEnOsFny8lUiOnTIoYL6cZl7h6xiaxmYpYjryQNtxs5S3x5LhoeZzEjyXC
qrcWoxmwnEER+qLkmTdxgcULoZceh2qrWw6/RpwCSUKlHZTEj5AmrbVS1t/qY3Wz
zCh+esjPLHQbeVJIfyd4sIsc/q1Aiip825/V69LfFD96K9DjbjHtwg025poZzsRz
X+zknOp4jkcQOu387xd24sSET/1rCB8jY7Y6P9WkNirpSM7bv4UDA9giTQIbP9Hb
`protect END_PROTECTED
