`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MG28XRBsjLKt2uCIPtAA/AjJRgg5aKz6Ok5jUafQY2U/1SQU7l35r9YGqcROu82/
nK8Ry1CgwYOx0gIdXWbgGiYbgnrMPm4hhPPReOLn/IrTax6LrUvZKVrYAUtwF0EZ
GlLp3duf8yoSX808VcyL/AIWa51s3vYwjzQZFmon1oUDEhvyR1mQXJmiFND1qV5R
cx0+Uz4yGr1ylkSyQv/sGg1U0XS56R9tbhO2cHFhh0m645XdVqhcAfdg5ovG2VKB
B+0oXx1VUwWH47+hLXz3VX0WUaHAxOKNwwcsWTelUePbKEeqKZLaL8IdzY9lU6D6
b6DgkY/50d82DtcMNc1ctNV0C3M4O5p0nlvwDhgLjBEv0MCKlNRCVb4JGjdX/99J
Ago/KfX2tISLFmJueL3G5CeNEO1aUrnEBwLLh9tP9f07dlyILLmpoUdpUZAIuJed
0FzOw0S/tjDwnG1Ut+JXGje7XtV0uQxgxvDWRLZZ0IKb3ZVp+gjow0BwgNM+E/dy
kUZ3ocpvK2J0ByUYfnmBOTmFpJSO6vZQxzCmXF3BuO9xnDkdr/7zsIXYc6mLzYCN
2YBg4UjMZSvL9O9OIzdblafBnGvNKpCxCRzyOODWous2vi7lJc0AqM+DKlc6qWh8
NhPnZJwNt+RdNTIYBT8Z0suV4KoY11wbK97TRzeRI31otSqapDtD82KjPfLdMrrM
CnvznHGKloT/C6Y0F+qiU6Nb1kwVy8I+GViQq09vlYsePN/6a+IiitMPW4vPtRrW
mBzNHOE1tHX1a0Ep89TMeNWbFDh7FwgUffazSP3baAe6GSMxffPFDfYFSUXNsSM5
E3+GJfHm3JPzgrDWevFI4XWFzYLBo4HKEPf8cZK5oACLjWnDn6pyp2VFCWOa48i/
NZPRXCXEZmzPer6M7YLdFuh7TzoOCswdjuStdJCxAtQUMbCvcTrkizNCkii6MGYU
aEtJrDwEKEKoFaeKBYt69dPap7jXWJKwpsMPt59iPZSQrf8fRBG8VhBTK8/ELY0n
R3X81IQvohw0ylEeV9+pd0CqafVOhC7hc6umKyzzGG16VVYQmBkrIx8QBduS7uuu
dL6wmAzZVlJcfZYAqdaKjLdHBfUE7GCa/Bhyt3ZUp8P20KtAj53qlw5bvFIXwmHf
x0BN1azHCuorwAFBUYxhZyCx5MuTTGgRKsReq7xnwhVcEEHIESWjMxYSE28ZTeVa
wsHevjqbZvor7FMCLDcU7Vz/feDXNMSSBqcxxSeuW4/b1CIO5VUlX0KihhMJMhWh
3NzQCNqC8xzdoee8vrhogIzJedeMH8Ib9PTIZWoglIk11rg9qttDGIo0pVkdXT5f
TpNd+sAhdcZB3VoejCNkwBz/T/xr/b/qv3qcUiwIqwSyHL42oSRTVJK3U7A02FeV
re1O1YbbndRHEcuu3Rc9CCYcHCTRoVUXaSMC55ckDHk4R9DVYXi6ZTCxfg5wYIhV
`protect END_PROTECTED
