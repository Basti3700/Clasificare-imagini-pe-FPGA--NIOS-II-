`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4WfStPdDBIZAC2+EPSRghtZWfrbDvlMwG7VhoI2r7UZYLc/d5//SZEe7tCjAyFwb
TUTGM9eVGDyK+kV/yJnWupDBafFuxAullMQCM1VKfrEU/FSlws+Ple0oxEEQS40N
UMyhCTXL74LBWpPYXBQi6T75EwwnHp7ClwuLt8rYrmcKgPKt1JT8T6zZJczsn5vX
9L0qx+8QVvN9dWzSS784u1m3K64wStBjWyfzpSVgm0ypx/7ndG0Oep7CQCk3M1Gt
8P2N2/iWXS6rgfwkYiJ3TxxD+RpYutfuFm8/yfCKy0kmo0/L6PSN7hxNHCPPqPcf
9WdCf4FHW9aASE2pp/KBa0Htkj5m4dpAj/3P+icYW0QE8OpN6FNRmS3ftKjqD6GC
Pkam2XHSw6DwRhbTQyIW48Za91C5S09EAItcdyEyuIH2q19X6CqWFO1u5xMBcFWT
WNUzgNrRFTgalBNKWsXC6P+ltjdCdPfPppz4tlssBCRa9B6UdabUFjQw58XH2Q8h
zAs28eypgWOYjPBXVWXR1uKuQkpZQ/3TeW8u5OqYWwgo7+v880Wc6VB6zC2ZgG9T
YVqPYWwmBUNkQINsRimeuSdG5QS2N3jSRphb2MAmF7T3EHYnk/6SPAelkOMUjQlK
4g2HOezefv7MVjZJxfTnRRhtEKxbcLCTWXsyO9R/Cfu2i5oAVbGvN3rWLJvAsNaY
t5OLKtb/UQUBKekZkVq5N3hPBVMQeILXLaEkfw/lulN/P0fiskDHjKlCrBlxbb51
PgfP5Pth12Ie904TQh3OccwTA5mqcCyXN6/OnKYSsp4bY6Dmj8n1PM3qpgdbcJt+
pChSPJfx4JkEDXKy0oNXJXUrb+DjV4ELoyvwLami1lTIUtsCx0Ei3ze2jDFsDdJP
13G49pEeHNQ6Jv/SUVqrYGSvH+q5K28s7O3HjeF4Qp483AuTredV/6If+FiYijRt
Og8dlGPhFETloIB/Bde22rDt9W2Zf1i7/W1tUljuqmOXUMY5Zw085HvF62isPoD4
2n1Kw0v5WwFywyjJdu9GRSj/qN4thxftbK2kZzv/1A/I1KoAWjMREC1Fbb5gnw2g
nx2OqvLAh2/tdmtwrx3Ll2jcFM3wler4XF31T/3Q6cGPwd4YVerupAw734Zg70ej
MWbXOGX1ULfARrYQBwnbz+T2cqdVZUAhzoRQ6Ik1MqwS04FwyZMG7/dPrInOCD9G
c6J9jw1JYfe6XuTvQVBwqcULXqTrPLThoNqN30LPZr4RI0LprI1dRPHxTR0Tepj6
oFc0GTHQRdVfIQp7o6fupay1PAvtfSXr+DacRub4hHxso74+qQd2UWqd2igV0/y+
nEFk5qnW4UT4ATy6mrkLCLdP1s8Frh6gjHZeijz2Tx6nzsBAb541/kcfJ4VG2U1v
inzzMfgybmCTJfm3Pylzvhb/yiJ/u4BMbQshCXvRXEhRP5PdXbWTBViIP9UILjZV
CLGY4bH97xwYHeWWeZsyq7Lme9HFxfb2b0z133AiMLqKlwZbai3A37Llr/wyM0Ei
XVEPGt5kz/G8zq0Cd6bPLQO3cfbosV2Y0WhvR0FAqv7tLc/DeEnMz820YXDOgbxf
q1IeY5GHrRqGp6K7fwyoGvaHhTFclNnWigYBLE+9kmb5qXdWMjGBP7IbsNG1gfHh
KB3j/mSYYm4wNFZ9cWP5j+HXDg0gdK/BKdHts7Wm6SakbTpUmd8/28vqP5kk82Dl
wLHi/bwm3x+uGKMDQRHXtzsPvb7sIXcopbnLACYwvETiI3P2x2P5/DtI7Ic786ww
KAdOe9jG+59l7sgpVXLn2/QH/yWUwxQLqqSSC6qRhBPtXayd8gcXMJ4eUE0Yw8aH
z94p9r2QOFy4S+IW2iLVic7pnWW22eNxOYSOpasEHFw6NsaV8fvtgvnjClT5O+FF
UtNYMi7rodbApARRN4CVLisZrOIB9S+UMOD87pQ0qXiMq8qVqD551MLJc2WZ9nrv
QGf3d9eKxDb7y4Q5lYBiOPn2znqry+/wSdzkNwlmetiogYJEd8raciF3Mn0tQc7u
te0PI+KeSZOeXaisCgzMoQKtTciQK5ZUWwbQrwaR0lpYudKBmmABhxHbPPINaszD
s2BpEWLEnsCVlj7z0AhGvXaSgnJ4Qd4X8Y5miPTSqZIU9D5SA6SR1f5BxVmvdT3T
aPKRO9HsBTIGIz5fio5tlhPsN+9eTPqyZx28yKKlLQKN/35pfaPStELoVJAJEyTR
3A6qDXT8dDaGmzZKZ55eFIn+qh2QDK/x+eXmYncD7etk3MsJ0L3rN17rPQkDRiAo
+QDmiKHow06NzjqWy5uD+yVdCYw85zgR/U21mZJsBI0=
`protect END_PROTECTED
