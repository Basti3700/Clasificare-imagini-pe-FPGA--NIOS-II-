library verilog;
use verilog.vl_types.all;
entity ama_coef_reg_ext_function is
    generic(
        width_coef      : integer := 1;
        register_clock_0: string  := "UNREGISTERED";
        register_aclr_0 : string  := "NONE";
        register_sclr_0 : string  := "NONE";
        register_clock_1: string  := "UNREGISTERED";
        register_aclr_1 : string  := "NONE";
        register_sclr_1 : string  := "NONE";
        register_clock_2: string  := "UNREGISTERED";
        register_aclr_2 : string  := "NONE";
        register_sclr_2 : string  := "NONE";
        register_clock_3: string  := "UNREGISTERED";
        register_aclr_3 : string  := "NONE";
        register_sclr_3 : string  := "NONE";
        number_of_multipliers: integer := 1;
        port_sign       : string  := "PORT_UNUSED";
        latency         : integer := 0;
        latency_clock_0 : string  := "UNREGISTERED";
        latency_aclr_0  : string  := "NONE";
        latency_sclr_0  : string  := "NONE";
        latency_clock_1 : string  := "UNREGISTERED";
        latency_aclr_1  : string  := "NONE";
        latency_sclr_1  : string  := "NONE";
        latency_clock_2 : string  := "UNREGISTERED";
        latency_aclr_2  : string  := "NONE";
        latency_sclr_2  : string  := "NONE";
        latency_clock_3 : string  := "UNREGISTERED";
        latency_aclr_3  : string  := "NONE";
        latency_sclr_3  : string  := "NONE";
        coef0_0         : vl_logic_vector;
        coef0_1         : vl_logic_vector;
        coef0_2         : vl_logic_vector;
        coef0_3         : vl_logic_vector;
        coef0_4         : vl_logic_vector;
        coef0_5         : vl_logic_vector;
        coef0_6         : vl_logic_vector;
        coef0_7         : vl_logic_vector;
        coef1_0         : vl_logic_vector;
        coef1_1         : vl_logic_vector;
        coef1_2         : vl_logic_vector;
        coef1_3         : vl_logic_vector;
        coef1_4         : vl_logic_vector;
        coef1_5         : vl_logic_vector;
        coef1_6         : vl_logic_vector;
        coef1_7         : vl_logic_vector;
        coef2_0         : vl_logic_vector;
        coef2_1         : vl_logic_vector;
        coef2_2         : vl_logic_vector;
        coef2_3         : vl_logic_vector;
        coef2_4         : vl_logic_vector;
        coef2_5         : vl_logic_vector;
        coef2_6         : vl_logic_vector;
        coef2_7         : vl_logic_vector;
        coef3_0         : vl_logic_vector;
        coef3_1         : vl_logic_vector;
        coef3_2         : vl_logic_vector;
        coef3_3         : vl_logic_vector;
        coef3_4         : vl_logic_vector;
        coef3_5         : vl_logic_vector;
        coef3_6         : vl_logic_vector;
        coef3_7         : vl_logic_vector
    );
    port(
        clock           : in     vl_logic_vector(3 downto 0);
        aclr            : in     vl_logic_vector(3 downto 0);
        sclr            : in     vl_logic_vector(3 downto 0);
        ena             : in     vl_logic_vector(3 downto 0);
        sign            : in     vl_logic;
        coefsel0        : in     vl_logic_vector(2 downto 0);
        coefsel1        : in     vl_logic_vector(2 downto 0);
        coefsel2        : in     vl_logic_vector(2 downto 0);
        coefsel3        : in     vl_logic_vector(2 downto 0);
        data_out_0      : out    vl_logic_vector;
        data_out_1      : out    vl_logic_vector;
        data_out_2      : out    vl_logic_vector;
        data_out_3      : out    vl_logic_vector
    );
    attribute coef0_0_mti_vect_attrib : integer;
    attribute coef0_0_mti_vect_attrib of coef0_0 : constant is 0;
    attribute coef0_1_mti_vect_attrib : integer;
    attribute coef0_1_mti_vect_attrib of coef0_1 : constant is 0;
    attribute coef0_2_mti_vect_attrib : integer;
    attribute coef0_2_mti_vect_attrib of coef0_2 : constant is 0;
    attribute coef0_3_mti_vect_attrib : integer;
    attribute coef0_3_mti_vect_attrib of coef0_3 : constant is 0;
    attribute coef0_4_mti_vect_attrib : integer;
    attribute coef0_4_mti_vect_attrib of coef0_4 : constant is 0;
    attribute coef0_5_mti_vect_attrib : integer;
    attribute coef0_5_mti_vect_attrib of coef0_5 : constant is 0;
    attribute coef0_6_mti_vect_attrib : integer;
    attribute coef0_6_mti_vect_attrib of coef0_6 : constant is 0;
    attribute coef0_7_mti_vect_attrib : integer;
    attribute coef0_7_mti_vect_attrib of coef0_7 : constant is 0;
    attribute coef1_0_mti_vect_attrib : integer;
    attribute coef1_0_mti_vect_attrib of coef1_0 : constant is 0;
    attribute coef1_1_mti_vect_attrib : integer;
    attribute coef1_1_mti_vect_attrib of coef1_1 : constant is 0;
    attribute coef1_2_mti_vect_attrib : integer;
    attribute coef1_2_mti_vect_attrib of coef1_2 : constant is 0;
    attribute coef1_3_mti_vect_attrib : integer;
    attribute coef1_3_mti_vect_attrib of coef1_3 : constant is 0;
    attribute coef1_4_mti_vect_attrib : integer;
    attribute coef1_4_mti_vect_attrib of coef1_4 : constant is 0;
    attribute coef1_5_mti_vect_attrib : integer;
    attribute coef1_5_mti_vect_attrib of coef1_5 : constant is 0;
    attribute coef1_6_mti_vect_attrib : integer;
    attribute coef1_6_mti_vect_attrib of coef1_6 : constant is 0;
    attribute coef1_7_mti_vect_attrib : integer;
    attribute coef1_7_mti_vect_attrib of coef1_7 : constant is 0;
    attribute coef2_0_mti_vect_attrib : integer;
    attribute coef2_0_mti_vect_attrib of coef2_0 : constant is 0;
    attribute coef2_1_mti_vect_attrib : integer;
    attribute coef2_1_mti_vect_attrib of coef2_1 : constant is 0;
    attribute coef2_2_mti_vect_attrib : integer;
    attribute coef2_2_mti_vect_attrib of coef2_2 : constant is 0;
    attribute coef2_3_mti_vect_attrib : integer;
    attribute coef2_3_mti_vect_attrib of coef2_3 : constant is 0;
    attribute coef2_4_mti_vect_attrib : integer;
    attribute coef2_4_mti_vect_attrib of coef2_4 : constant is 0;
    attribute coef2_5_mti_vect_attrib : integer;
    attribute coef2_5_mti_vect_attrib of coef2_5 : constant is 0;
    attribute coef2_6_mti_vect_attrib : integer;
    attribute coef2_6_mti_vect_attrib of coef2_6 : constant is 0;
    attribute coef2_7_mti_vect_attrib : integer;
    attribute coef2_7_mti_vect_attrib of coef2_7 : constant is 0;
    attribute coef3_0_mti_vect_attrib : integer;
    attribute coef3_0_mti_vect_attrib of coef3_0 : constant is 0;
    attribute coef3_1_mti_vect_attrib : integer;
    attribute coef3_1_mti_vect_attrib of coef3_1 : constant is 0;
    attribute coef3_2_mti_vect_attrib : integer;
    attribute coef3_2_mti_vect_attrib of coef3_2 : constant is 0;
    attribute coef3_3_mti_vect_attrib : integer;
    attribute coef3_3_mti_vect_attrib of coef3_3 : constant is 0;
    attribute coef3_4_mti_vect_attrib : integer;
    attribute coef3_4_mti_vect_attrib of coef3_4 : constant is 0;
    attribute coef3_5_mti_vect_attrib : integer;
    attribute coef3_5_mti_vect_attrib of coef3_5 : constant is 0;
    attribute coef3_6_mti_vect_attrib : integer;
    attribute coef3_6_mti_vect_attrib of coef3_6 : constant is 0;
    attribute coef3_7_mti_vect_attrib : integer;
    attribute coef3_7_mti_vect_attrib of coef3_7 : constant is 0;
end ama_coef_reg_ext_function;
